`default_nettype none
/*
 *  SPDX-FileCopyrightText: 2017 Clifford Wolf
 *
 *  PicoSoC - A simple example SoC using PicoRV32
 *
 *  Copyright (C) 2017  Clifford Wolf <clifford@clifford.at>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 *  SPDX-License-Identifier: ISC
 */

`timescale 1 ns / 1 ps

/* tbuart --- mimic an external UART display, operating at 9600 baud	*/
/* and accepting ASCII characters for display.				*/

/* To do:  Match a known UART 3.3V 16x2 LCD display.  However, it	*/
/* should be possible on a testing system to interface to the UART	*/
/* pins on a Raspberry Pi, also running at 3.3V.			*/

module tbuart (
	input  ser_rx,
	output  ser_tx
);
	reg [3:0] recv_state;
	reg [2:0] recv_divcnt;
	reg [7:0] recv_pattern;
	reg [8*50-1:0] recv_buf_data;	// 50 characters.  Increase as needed for tests.

	reg clk;

	initial begin
		clk <= 1'b0;
		recv_state <= 0;
		recv_divcnt <= 0;
		recv_pattern <= 0;
		recv_buf_data <= 0;
	end

	// NOTE:  Running at 3.0us clock period @ 5 clocks per bit = 15.0us per
	// bit ~= 64 kbaud. Not tuned to any particular UART.  Most run at
	// 9600 baud default and will bounce up to higher baud rates when
	// passed specific command words.

//	always #1500 clk <= (clk === 1'b0);
	always #2650 clk <= (clk === 1'b0);  // working for 9600 baud
//	always #125 clk <= (clk === 1'b0);

	always @(posedge clk) begin
		recv_divcnt <= recv_divcnt + 1;
		case (recv_state)
			0: begin
				if (!ser_rx)
					recv_state <= 1;
				recv_divcnt <= 0;
			end
			1: begin
				if (2*recv_divcnt > 3'd3) begin
					recv_state <= 2;
					recv_divcnt <= 0;
				end
			end
			10: begin
				if (recv_divcnt > 3'd3) begin
					// 0x0a = '\n'
					if (recv_pattern == 8'h0a) begin
						$display("output: %s", recv_buf_data);
					end else begin
						recv_buf_data <= {recv_buf_data, recv_pattern};
					end
					recv_state <= 0;
				end
			end
			default: begin
				if (recv_divcnt > 3'd3) begin
					recv_pattern <= {ser_rx, recv_pattern[7:1]};
					recv_state <= recv_state + 1;
					recv_divcnt <= 0;
				end
			end
		endcase
	end

endmodule
`default_nettype none
/*
 *  SPDX-FileCopyrightText: 2017 Clifford Wolf
 *
 *  PicoSoC - A simple example SoC using PicoRV32
 *
 *  Copyright (C) 2017  Clifford Wolf <clifford@clifford.at>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 *  SPDX-License-Identifier: ISC
 */

`timescale 1 ns / 1 ps

//
// Simple SPI flash simulation model
//
// This model samples io input signals 1ns before the SPI clock edge and
// updates output signals 1ns after the SPI clock edge.
//
// Supported commands:
//    AB, B9, FF, 03, BB, EB, ED
//
// Well written SPI flash data sheets:
//    Cypress S25FL064L http://www.cypress.com/file/316661/download
//    Cypress S25FL128L http://www.cypress.com/file/316171/download
//

module spiflash #(
	parameter FILENAME = "firmware.hex"
)(
	input csb,
	input clk,
	inout io0, // MOSI
	inout io1, // MISO
	inout io2,
	inout io3
);
	localparam verbose = 0;
	localparam integer latency = 8;
	
	reg [7:0] buffer;
	reg [3:0] reset_count = 0;
	reg [3:0] reset_monitor = 0;
	integer bitcount = 0;
	integer bytecount = 0;
	integer dummycount = 0;

	reg [7:0] spi_cmd;
	reg [7:0] xip_cmd = 0;
	reg [23:0] spi_addr;

	reg [7:0] spi_in;
	reg [7:0] spi_out;
	reg spi_io_vld;

	reg powered_up = 1;

	localparam [3:0] mode_spi         = 1;
	localparam [3:0] mode_dspi_rd     = 2;
	localparam [3:0] mode_dspi_wr     = 3;
	localparam [3:0] mode_qspi_rd     = 4;
	localparam [3:0] mode_qspi_wr     = 5;
	localparam [3:0] mode_qspi_ddr_rd = 6;
	localparam [3:0] mode_qspi_ddr_wr = 7;

	reg [3:0] mode = 0;
	reg [3:0] next_mode = 0;

	reg io0_oe = 0;
	reg io1_oe = 0;
	reg io2_oe = 0;
	reg io3_oe = 0;

	reg io0_dout = 0;
	reg io1_dout = 0;
	reg io2_dout = 0;
	reg io3_dout = 0;

	assign #1 io0 = io0_oe ? io0_dout : 1'bz;
	assign #1 io1 = io1_oe ? io1_dout : 1'bz;
	assign #1 io2 = io2_oe ? io2_dout : 1'bz;
	assign #1 io3 = io3_oe ? io3_dout : 1'bz;

	wire io0_delayed;
	wire io1_delayed;
	wire io2_delayed;
	wire io3_delayed;

	assign #1 io0_delayed = io0;
	assign #1 io1_delayed = io1;
	assign #1 io2_delayed = io2;
	assign #1 io3_delayed = io3;

	// 16 MB (128Mb) Flash
	reg [7:0] memory [0:16*1024*1024-1];

	initial begin
		$display("Reading %s",  FILENAME);
		$readmemh(FILENAME, memory);
		//$display("Memory 5 bytes = 0x%02x 0x%02x 0x%02x 0x%02x 0x%02x",
		//	memory[0], memory[1], memory[2],
		//	memory[3], memory[4]);
		$display("%s loaded into memory", FILENAME);
		$display("Memory 5 bytes = 0x%02x 0x%02x 0x%02x 0x%02x 0x%02x",
			memory[0], memory[1], memory[2],
			memory[3], memory[4]);
	end

	task spi_action;
		begin
			spi_in = buffer;

			if (bytecount == 1) begin
				spi_cmd = buffer;

				if (spi_cmd == 8'h ab)
					powered_up = 1;

				if (spi_cmd == 8'h b9)
					powered_up = 0;

				if (spi_cmd == 8'h ff)
					xip_cmd = 0;
			end

			if (powered_up && spi_cmd == 'h 03) begin
				if (bytecount == 2)
					spi_addr[23:16] = buffer;

				if (bytecount == 3)
					spi_addr[15:8] = buffer;

				if (bytecount == 4)
					spi_addr[7:0] = buffer;

				if (bytecount >= 4) begin
					buffer = memory[spi_addr];
					spi_addr = spi_addr + 1;
				end
			end

			if (powered_up && spi_cmd == 'h bb) begin
				if (bytecount == 1)
					mode = mode_dspi_rd;

				if (bytecount == 2)
					spi_addr[23:16] = buffer;

				if (bytecount == 3)
					spi_addr[15:8] = buffer;

				if (bytecount == 4)
					spi_addr[7:0] = buffer;

				if (bytecount == 5) begin
					xip_cmd = (buffer == 8'h a5) ? spi_cmd : 8'h 00;
					mode = mode_dspi_wr;
					dummycount = latency;
				end

				if (bytecount >= 5) begin
					buffer = memory[spi_addr];
					spi_addr = spi_addr + 1;
				end
			end

			if (powered_up && spi_cmd == 'h eb) begin
				if (bytecount == 1)
					mode = mode_qspi_rd;

				if (bytecount == 2)
					spi_addr[23:16] = buffer;

				if (bytecount == 3)
					spi_addr[15:8] = buffer;

				if (bytecount == 4)
					spi_addr[7:0] = buffer;

				if (bytecount == 5) begin
					xip_cmd = (buffer == 8'h a5) ? spi_cmd : 8'h 00;
					mode = mode_qspi_wr;
					dummycount = latency;
				end

				if (bytecount >= 5) begin
					buffer = memory[spi_addr];
					spi_addr = spi_addr + 1;
				end
			end

			if (powered_up && spi_cmd == 'h ed) begin
				if (bytecount == 1)
					next_mode = mode_qspi_ddr_rd;

				if (bytecount == 2)
					spi_addr[23:16] = buffer;

				if (bytecount == 3)
					spi_addr[15:8] = buffer;

				if (bytecount == 4)
					spi_addr[7:0] = buffer;

				if (bytecount == 5) begin
					xip_cmd = (buffer == 8'h a5) ? spi_cmd : 8'h 00;
					mode = mode_qspi_ddr_wr;
					dummycount = latency;
				end

				if (bytecount >= 5) begin
					buffer = memory[spi_addr];
					spi_addr = spi_addr + 1;
				end
			end

			spi_out = buffer;
			spi_io_vld = 1;

			if (verbose) begin
				if (bytecount == 1)
					$write("<SPI-START>");
				$write("<SPI:%02x:%02x>", spi_in, spi_out);
			end

		end
	endtask

	task ddr_rd_edge;
		begin
			buffer = {buffer, io3_delayed, io2_delayed, io1_delayed, io0_delayed};
			bitcount = bitcount + 4;
			if (bitcount == 8) begin
				bitcount = 0;
				bytecount = bytecount + 1;
				spi_action;
			end
		end
	endtask

	task ddr_wr_edge;
		begin
			io0_oe = 1;
			io1_oe = 1;
			io2_oe = 1;
			io3_oe = 1;

			io0_dout = buffer[4];
			io1_dout = buffer[5];
			io2_dout = buffer[6];
			io3_dout = buffer[7];

			buffer = {buffer, 4'h 0};
			bitcount = bitcount + 4;
			if (bitcount == 8) begin
				bitcount = 0;
				bytecount = bytecount + 1;
				spi_action;
			end
		end
	endtask

	always @(csb) begin
		if (csb) begin
			if (verbose) begin
				$display("");
				$fflush;
			end
			buffer = 0;
			bitcount = 0;
			bytecount = 0;
			mode = mode_spi;
			io0_oe = 0;
			io1_oe = 0;
			io2_oe = 0;
			io3_oe = 0;

			// Handle MBR.  If in XIP continuous mode, the following
			// 8 clock cycles are normally not expected to be a command.
			// If followed by CSB high, however, if the address bits
			// are consistent with io0 == 1 for 8 clk cycles, then an
			// MBR has been issued and the system must exit XIP
			// continuous mode.
			if (xip_cmd == 8'hbb || xip_cmd == 8'heb
					|| xip_cmd == 8'hed) begin
				if (reset_count == 4'h8 && reset_monitor == 4'h8) begin
					xip_cmd = 8'h00;
					spi_cmd = 8'h03;
				end
			end
		end else
		if (xip_cmd) begin
			buffer = xip_cmd;
			bitcount = 0;
			bytecount = 1;
			spi_action;
		end
	end

	always @(posedge clk or posedge csb) begin
		if (csb == 1'b1) begin
			reset_count = 0;
			reset_monitor = 0;
		end else begin
			if (reset_count < 4'h9) begin
				reset_count = reset_count + 1;
				if (io0_delayed == 1'b1) begin
				    reset_monitor = reset_monitor + 1;
				end
			end
		end
	end

	always @(csb, clk) begin
		spi_io_vld = 0;
		if (!csb && !clk) begin
			if (dummycount > 0) begin
				io0_oe = 0;
				io1_oe = 0;
				io2_oe = 0;
				io3_oe = 0;
			end else
			case (mode)
				mode_spi: begin
					io0_oe = 0;
					io1_oe = 1;
					io2_oe = 0;
					io3_oe = 0;
					io1_dout = buffer[7];
				end
				mode_dspi_rd: begin
					io0_oe = 0;
					io1_oe = 0;
					io2_oe = 0;
					io3_oe = 0;
				end
				mode_dspi_wr: begin
					io0_oe = 1;
					io1_oe = 1;
					io2_oe = 0;
					io3_oe = 0;
					io0_dout = buffer[6];
					io1_dout = buffer[7];
				end
				mode_qspi_rd: begin
					io0_oe = 0;
					io1_oe = 0;
					io2_oe = 0;
					io3_oe = 0;
				end
				mode_qspi_wr: begin
					io0_oe = 1;
					io1_oe = 1;
					io2_oe = 1;
					io3_oe = 1;
					io0_dout = buffer[4];
					io1_dout = buffer[5];
					io2_dout = buffer[6];
					io3_dout = buffer[7];
				end
				mode_qspi_ddr_rd: begin
					ddr_rd_edge;
				end
				mode_qspi_ddr_wr: begin
					ddr_wr_edge;
				end
			endcase
			if (next_mode) begin
				case (next_mode)
					mode_qspi_ddr_rd: begin
						io0_oe = 0;
						io1_oe = 0;
						io2_oe = 0;
						io3_oe = 0;
					end
					mode_qspi_ddr_wr: begin
						io0_oe = 1;
						io1_oe = 1;
						io2_oe = 1;
						io3_oe = 1;
						io0_dout = buffer[4];
						io1_dout = buffer[5];
						io2_dout = buffer[6];
						io3_dout = buffer[7];
					end
				endcase
				mode = next_mode;
				next_mode = 0;
			end
		end
	end

	always @(posedge clk) begin
		if (!csb) begin
			if (dummycount > 0) begin
				dummycount = dummycount - 1;
			end else
			case (mode)
				mode_spi: begin
					buffer = {buffer, io0};
					bitcount = bitcount + 1;
					if (bitcount == 8) begin
						bitcount = 0;
						bytecount = bytecount + 1;
						spi_action;
					end
				end
				mode_dspi_rd, mode_dspi_wr: begin
					buffer = {buffer, io1, io0};
					bitcount = bitcount + 2;
					if (bitcount == 8) begin
						bitcount = 0;
						bytecount = bytecount + 1;
						spi_action;
					end
				end
				mode_qspi_rd, mode_qspi_wr: begin
					buffer = {buffer, io3, io2, io1, io0};
					bitcount = bitcount + 4;
					if (bitcount == 8) begin
						bitcount = 0;
						bytecount = bytecount + 1;
						spi_action;
					end
				end
				mode_qspi_ddr_rd: begin
					ddr_rd_edge;
				end
				mode_qspi_ddr_wr: begin
					ddr_wr_edge;
				end
			endcase
		end
	end
endmodule
`default_nettype none

`timescale 1 ns / 1 ps

module wb_rw_test(
    input wire rx,
    output wire tx,
    input wire start
);

//parameter BTIME = 8680;
parameter BTIME = 2175;
//parameter BTIME = 2177;
reg TX;
wire RX;

reg [31:0] data;

assign RX = rx;
assign tx = TX;

initial begin
    TX <= 1'b1;
    #10000;
    $display("Executing SRAM write");
    wb_write(30'h00400024, 32'h775555ab);
    $display("Executing SRAM read");
    wb_read (32'h00400024, data);
    $display("output: %h", data);

    if (data != 32'h775555ab) begin
        $display("SRAM write failed");
        $finish;
    end else begin
        $display("SRAM write succeeded");
    end
end

task uart_put(input [7:0] b);
    integer i;
    begin
        TX = 1'b0;
        #BTIME;
        for(i=0; i<8; i=i+1) begin
            TX = b[i];
            #BTIME;
        end
        TX = 1'b1;
        #(BTIME);
    end
endtask

task uart_put_ns(input [7:0] b);
    integer i;
    begin
        TX = 1'b0;
        #BTIME;
        for(i=0; i<8; i=i+1) begin
            TX = b[i];
            #BTIME;
        end
        TX = 1'b1;
//        #(BTIME);
    end
endtask

task uart_get(output [7:0] b);
    integer i;
    begin
        @(negedge RX);
        #BTIME;
        for(i=0; i<8; i=i+1) begin
            #(BTIME/2);
            b[i] <= RX;
            #(BTIME/2);
        end
        #(BTIME);
    end
endtask

task wb_read (input [31:0] addr, output [31:0] word);
    begin
        uart_put(8'h2);     // read cmd
        uart_put(8'h1);      // size
        uart_put(addr[31:24]);
        uart_put(addr[23:16]);
        uart_put(addr[15:8]);
        uart_put_ns(addr[7:0]);
        uart_get(word[31:24]);
        uart_get(word[23:16]);
        uart_get(word[15:8]);
        uart_get(word[7:0]);
    end
endtask

task wb_write (input [31:0] addr, input [31:0] word);
    begin
        uart_put(8'h1);     // write cmd
        uart_put(8'h1);      // size
        uart_put(addr[31:24]);
        uart_put(addr[23:16]);
        uart_put(addr[15:8]);
        uart_put(addr[7:0]);
        uart_put(word[31:24]);
        uart_put(word[23:16]);
        uart_put(word[15:8]);
        uart_put(word[7:0]);
    end
endtask

endmodule
module RAM256 #( parameter COLS=1)
(

    VPWR,
    VGND,

    CLK,
    WE0,
    EN0,
    Di0,
    Do0,
    A0
);
    localparam A_WIDTH = 8+$clog2(COLS);

    input   wire            VPWR;
    input   wire            VGND;
    input   wire            CLK;
    input   wire    [3:0]   WE0;
    input   wire            EN0;
    input   wire    [31:0]  Di0;
    output  reg     [31:0]  Do0;
    input   wire    [(A_WIDTH - 1): 0]   A0;

    reg [31:0] RAM[(256*COLS)-1 : 0];

    always @(posedge CLK)
        if(EN0) begin
            Do0 <= RAM[A0];
            if(WE0[0]) RAM[A0][ 7: 0] <= Di0[7:0];
            if(WE0[1]) RAM[A0][15:8] <= Di0[15:8];
            if(WE0[2]) RAM[A0][23:16] <= Di0[23:16];
            if(WE0[3]) RAM[A0][31:24] <= Di0[31:24];
        end
        else
            Do0 <= 32'b0;

endmodule
module RAM128 #( parameter COLS=1)
(

    VPWR,
    VGND,

    CLK,
    WE0,
    EN0,
    Di0,
    Do0,
    A0
);
    localparam A_WIDTH = 7+$clog2(COLS);

    input   wire            VPWR;
    input   wire            VGND;
    input   wire            CLK;
    input   wire    [3:0]   WE0;
    input   wire            EN0;
    input   wire    [31:0]  Di0;
    output  reg     [31:0]  Do0;
    input   wire    [(A_WIDTH - 1): 0]   A0;

    reg [31:0] RAM[(256*COLS)-1 : 0];

    always @(posedge CLK)
        if(EN0) begin
            Do0 <= RAM[A0];
            if(WE0[0]) RAM[A0][ 7: 0] <= Di0[7:0];
            if(WE0[1]) RAM[A0][15:8] <= Di0[15:8];
            if(WE0[2]) RAM[A0][23:16] <= Di0[23:16];
            if(WE0[3]) RAM[A0][31:24] <= Di0[31:24];
        end
        else
            Do0 <= 32'b0;

endmodule
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0



// Global parameters










// Analog pads are only used by the "caravan" module and associated
// modules such as user_analog_project_wrapper and chip_io_alt.






// Size of soc_mem_synth

// Type and size of soc_mem
// `define USE_OPENRAM

// don't change the following without double checking addr widths


// Number of columns in the custom memory; takes one of three values:
// 1 column : 1 KB, 2 column: 2 KB, 4 column: 4KB



// not really parameterized but just to easily keep track of the number
// of ram_block across different modules


// Clock divisor default value


// GPIO control default mode and enable for most I/Os
// Most I/Os set to be user bidirectional pins on power-up.











 // __GLOBAL_DEFINE_H
//--------------------------------------------------------------------------------
// Auto-generated by Migen (9a0be7a) & LiteX (470fc6f) on 2022-10-14 12:53:55
//--------------------------------------------------------------------------------
module mgmt_core(

    inout VPWR,	    /* 1.8V domain */
    inout VGND,

	input wire core_clk,
	input wire core_rstn,
	output wire flash_cs_n,
	output reg flash_clk,
	output reg flash_io0_oeb,
	output wire flash_io1_oeb,
	output wire flash_io2_oeb,
	output wire flash_io3_oeb,
	output reg flash_io0_do,
	output wire flash_io1_do,
	output wire flash_io2_do,
	output wire flash_io3_do,
	input wire flash_io0_di,
	input wire flash_io1_di,
	input wire flash_io2_di,
	input wire flash_io3_di,
	output reg spi_clk,
	output reg spi_cs_n,
	output reg spi_mosi,
	input wire spi_miso,
	output wire spi_sdoenb,
	output wire mprj_wb_iena,
	output wire mprj_cyc_o,
	output wire mprj_stb_o,
	output wire mprj_we_o,
	output wire [3:0] mprj_sel_o,
	output reg [31:0] mprj_adr_o,
	output wire [31:0] mprj_dat_o,
	input wire [31:0] mprj_dat_i,
	input wire mprj_ack_i,
	input wire [31:0] hk_dat_i,
	output wire hk_stb_o,
	output wire hk_cyc_o,
	input wire hk_ack_i,
	output reg serial_tx,
	input wire serial_rx,
	input wire debug_in,
	output wire debug_out,
	output wire debug_oeb,
	output wire debug_mode,
	output wire uart_enabled,
	output wire gpio_out_pad,
	input wire gpio_in_pad,
	output wire gpio_outenb_pad,
	output wire gpio_inenb_pad,
	output wire gpio_mode0_pad,
	output wire gpio_mode1_pad,
	output reg [127:0] la_output,
	input wire [127:0] la_input,
	output reg [127:0] la_oenb,
	output reg [127:0] la_iena,
	output wire qspi_enabled,
	output wire spi_enabled,
	output wire trap,
	output wire [2:0] user_irq_ena,
	input wire [5:0] user_irq,
	input wire clk_in,
	output wire clk_out,
	input wire resetn_in,
	output wire resetn_out,
	input wire serial_load_in,
	output wire serial_load_out,
	input wire serial_data_2_in,
	output wire serial_data_2_out,
	input wire serial_resetn_in,
	output wire serial_resetn_out,
	input wire serial_clock_in,
	output wire serial_clock_out,
	input wire rstb_l_in,
	output wire rstb_l_out,
	input wire por_l_in,
	output wire por_l_out,
	input wire porb_h_in,
	output wire porb_h_out
);

wire core_rst;
wire sys_clk;
wire sys_rst;
wire por_clk;
reg int_rst = 1'd1;
reg mgmtsoc_soc_rst = 1'd0;
wire mgmtsoc_cpu_rst;
reg [1:0] mgmtsoc_reset_storage = 2'd0;
reg mgmtsoc_reset_re = 1'd0;
reg [31:0] mgmtsoc_scratch_storage = 32'd305419896;
reg mgmtsoc_scratch_re = 1'd0;
wire [31:0] mgmtsoc_bus_errors_status;
wire mgmtsoc_bus_errors_we;
reg mgmtsoc_bus_errors_re = 1'd0;
wire mgmtsoc_bus_error;
reg [31:0] mgmtsoc_bus_errors = 32'd0;
wire mgmtsoc_reset;
reg [31:0] mgmtsoc_interrupt = 32'd0;
wire [29:0] mgmtsoc_ibus_ibus_adr;
wire [31:0] mgmtsoc_ibus_ibus_dat_w;
wire [31:0] mgmtsoc_ibus_ibus_dat_r;
wire [3:0] mgmtsoc_ibus_ibus_sel;
wire mgmtsoc_ibus_ibus_cyc;
wire mgmtsoc_ibus_ibus_stb;
wire mgmtsoc_ibus_ibus_ack;
wire mgmtsoc_ibus_ibus_we;
wire [2:0] mgmtsoc_ibus_ibus_cti;
wire [1:0] mgmtsoc_ibus_ibus_bte;
wire mgmtsoc_ibus_ibus_err;
wire [29:0] mgmtsoc_dbus_dbus_adr;
wire [31:0] mgmtsoc_dbus_dbus_dat_w;
wire [31:0] mgmtsoc_dbus_dbus_dat_r;
wire [3:0] mgmtsoc_dbus_dbus_sel;
wire mgmtsoc_dbus_dbus_cyc;
wire mgmtsoc_dbus_dbus_stb;
wire mgmtsoc_dbus_dbus_ack;
wire mgmtsoc_dbus_dbus_we;
wire [2:0] mgmtsoc_dbus_dbus_cti;
wire [1:0] mgmtsoc_dbus_dbus_bte;
wire mgmtsoc_dbus_dbus_err;
reg mgmtsoc_vexriscv_debug_reset = 1'd0;
reg mgmtsoc_vexriscv_ibus_err = 1'd0;
reg mgmtsoc_vexriscv_dbus_err = 1'd0;
reg mgmtsoc_vexriscv_i_cmd_valid = 1'd0;
reg mgmtsoc_vexriscv_i_cmd_payload_wr = 1'd0;
reg [7:0] mgmtsoc_vexriscv_i_cmd_payload_address = 8'd0;
reg [31:0] mgmtsoc_vexriscv_i_cmd_payload_data = 32'd0;
wire mgmtsoc_vexriscv_o_cmd_ready;
wire [31:0] mgmtsoc_vexriscv_o_rsp_data;
wire mgmtsoc_vexriscv_o_resetOut;
reg mgmtsoc_vexriscv_reset_debug_logic = 1'd0;
reg mgmtsoc_vexriscv_transfer_complete = 1'd0;
reg mgmtsoc_vexriscv_transfer_in_progress = 1'd0;
reg mgmtsoc_vexriscv_transfer_wait_for_ack = 1'd0;
wire [29:0] mgmtsoc_vexriscv_debug_bus_adr;
wire [31:0] mgmtsoc_vexriscv_debug_bus_dat_w;
reg [31:0] mgmtsoc_vexriscv_debug_bus_dat_r = 32'd0;
wire [3:0] mgmtsoc_vexriscv_debug_bus_sel;
wire mgmtsoc_vexriscv_debug_bus_cyc;
wire mgmtsoc_vexriscv_debug_bus_stb;
reg mgmtsoc_vexriscv_debug_bus_ack = 1'd0;
wire mgmtsoc_vexriscv_debug_bus_we;
wire [2:0] mgmtsoc_vexriscv_debug_bus_cti;
wire [1:0] mgmtsoc_vexriscv_debug_bus_bte;
reg mgmtsoc_vexriscv_debug_bus_err = 1'd0;
reg [31:0] mgmtsoc_vexriscv = 32'd268435456;
reg [31:0] mgmtsoc_load_storage = 32'd0;
reg mgmtsoc_load_re = 1'd0;
reg [31:0] mgmtsoc_reload_storage = 32'd0;
reg mgmtsoc_reload_re = 1'd0;
reg mgmtsoc_en_storage = 1'd0;
reg mgmtsoc_en_re = 1'd0;
reg mgmtsoc_update_value_storage = 1'd0;
reg mgmtsoc_update_value_re = 1'd0;
reg [31:0] mgmtsoc_value_status = 32'd0;
wire mgmtsoc_value_we;
reg mgmtsoc_value_re = 1'd0;
wire mgmtsoc_irq;
wire mgmtsoc_zero_status;
reg mgmtsoc_zero_pending = 1'd0;
wire mgmtsoc_zero_trigger;
reg mgmtsoc_zero_clear = 1'd0;
reg mgmtsoc_zero_trigger_d = 1'd0;
wire mgmtsoc_zero0;
wire mgmtsoc_status_status;
wire mgmtsoc_status_we;
reg mgmtsoc_status_re = 1'd0;
wire mgmtsoc_zero1;
wire mgmtsoc_pending_status;
wire mgmtsoc_pending_we;
reg mgmtsoc_pending_re = 1'd0;
reg mgmtsoc_pending_r = 1'd0;
wire mgmtsoc_zero2;
reg mgmtsoc_enable_storage = 1'd0;
reg mgmtsoc_enable_re = 1'd0;
reg [31:0] mgmtsoc_value = 32'd0;
wire [29:0] dff_bus_adr;
wire [31:0] dff_bus_dat_w;
wire [31:0] dff_bus_dat_r;
wire [3:0] dff_bus_sel;
wire dff_bus_cyc;
wire dff_bus_stb;
reg dff_bus_ack = 1'd0;
wire dff_bus_we;
wire [2:0] dff_bus_cti;
wire [1:0] dff_bus_bte;
reg dff_bus_err = 1'd0;
wire [31:0] dff_di;
wire [31:0] dff_do;
reg [3:0] dff_we = 4'd0;
wire dff_en;
wire [29:0] dff2_bus_adr;
wire [31:0] dff2_bus_dat_w;
wire [31:0] dff2_bus_dat_r;
wire [3:0] dff2_bus_sel;
wire dff2_bus_cyc;
wire dff2_bus_stb;
reg dff2_bus_ack = 1'd0;
wire dff2_bus_we;
wire [2:0] dff2_bus_cti;
wire [1:0] dff2_bus_bte;
reg dff2_bus_err = 1'd0;
wire [31:0] dff2_di;
wire [31:0] dff2_do;
reg [3:0] dff2_we = 4'd0;
wire dff2_en;
reg mgmtsoc_litespisdrphycore_source_valid = 1'd0;
wire mgmtsoc_litespisdrphycore_source_ready;
reg mgmtsoc_litespisdrphycore_source_first = 1'd0;
reg mgmtsoc_litespisdrphycore_source_last = 1'd0;
wire [31:0] mgmtsoc_litespisdrphycore_source_payload_data;
wire mgmtsoc_litespisdrphycore_sink_valid;
reg mgmtsoc_litespisdrphycore_sink_ready = 1'd0;
wire mgmtsoc_litespisdrphycore_sink_first;
wire mgmtsoc_litespisdrphycore_sink_last;
wire [31:0] mgmtsoc_litespisdrphycore_sink_payload_data;
wire [5:0] mgmtsoc_litespisdrphycore_sink_payload_len;
wire [3:0] mgmtsoc_litespisdrphycore_sink_payload_width;
wire [7:0] mgmtsoc_litespisdrphycore_sink_payload_mask;
wire mgmtsoc_litespisdrphycore_cs;
wire [7:0] mgmtsoc_litespisdrphycore_spi_clk_divisor;
reg [7:0] mgmtsoc_litespisdrphycore_storage = 8'd1;
reg mgmtsoc_litespisdrphycore_re = 1'd0;
wire [7:0] mgmtsoc_litespisdrphycore_div;
wire [7:0] mgmtsoc_litespisdrphycore_sample_cnt;
wire [7:0] mgmtsoc_litespisdrphycore_update_cnt;
wire mgmtsoc_litespisdrphycore_posedge;
wire mgmtsoc_litespisdrphycore_negedge;
wire mgmtsoc_litespisdrphycore_sample;
wire mgmtsoc_litespisdrphycore_update;
reg mgmtsoc_litespisdrphycore_en = 1'd0;
reg [7:0] mgmtsoc_litespisdrphycore_cnt = 8'd0;
reg mgmtsoc_litespisdrphycore_en_int = 1'd0;
reg mgmtsoc_litespisdrphycore_clk = 1'd0;
reg mgmtsoc_litespisdrphycore_posedge_reg = 1'd0;
reg mgmtsoc_litespisdrphycore_posedge_reg2 = 1'd0;
wire mgmtsoc_litespisdrphycore_wait;
wire mgmtsoc_litespisdrphycore_done;
reg [3:0] mgmtsoc_litespisdrphycore_count = 4'd11;
wire mgmtsoc_litespisdrphycore_cs_enable;
reg mgmtsoc_litespisdrphycore_dq_o = 1'd0;
reg [1:0] mgmtsoc_litespisdrphycore_dq_i = 2'd0;
wire mgmtsoc_litespisdrphycore_dq_oe;
reg [7:0] mgmtsoc_litespisdrphycore_sr_cnt = 8'd0;
reg mgmtsoc_litespisdrphycore_sr_out_load = 1'd0;
reg mgmtsoc_litespisdrphycore_sr_out_shift = 1'd0;
reg [31:0] mgmtsoc_litespisdrphycore_sr_out = 32'd0;
reg mgmtsoc_litespisdrphycore_sr_in_shift = 1'd0;
reg [31:0] mgmtsoc_litespisdrphycore_sr_in = 32'd0;
reg mgmtsoc_litespisdrphycore0 = 1'd0;
reg [1:0] mgmtsoc_litespisdrphycore1 = 2'd0;
reg [3:0] mgmtsoc_litespisdrphycore2 = 4'd0;
reg [7:0] mgmtsoc_litespisdrphycore3 = 8'd0;
wire mgmtsoc_crossbar_source_valid;
wire mgmtsoc_crossbar_source_ready;
wire mgmtsoc_crossbar_source_first;
wire mgmtsoc_crossbar_source_last;
wire [31:0] mgmtsoc_crossbar_source_payload_data;
wire [5:0] mgmtsoc_crossbar_source_payload_len;
wire [3:0] mgmtsoc_crossbar_source_payload_width;
wire [7:0] mgmtsoc_crossbar_source_payload_mask;
wire mgmtsoc_crossbar_sink_valid;
wire mgmtsoc_crossbar_sink_ready;
wire mgmtsoc_crossbar_sink_first;
wire mgmtsoc_crossbar_sink_last;
wire [31:0] mgmtsoc_crossbar_sink_payload_data;
reg mgmtsoc_crossbar_cs = 1'd0;
reg mgmtsoc_litespimmap_source_valid = 1'd0;
wire mgmtsoc_litespimmap_source_ready;
reg mgmtsoc_litespimmap_source_first = 1'd0;
reg mgmtsoc_litespimmap_source_last = 1'd0;
reg [31:0] mgmtsoc_litespimmap_source_payload_data = 32'd0;
reg [5:0] mgmtsoc_litespimmap_source_payload_len = 6'd0;
reg [3:0] mgmtsoc_litespimmap_source_payload_width = 4'd0;
reg [7:0] mgmtsoc_litespimmap_source_payload_mask = 8'd0;
wire mgmtsoc_litespimmap_sink_valid;
reg mgmtsoc_litespimmap_sink_ready = 1'd0;
wire mgmtsoc_litespimmap_sink_first;
wire mgmtsoc_litespimmap_sink_last;
wire [31:0] mgmtsoc_litespimmap_sink_payload_data;
wire [29:0] mgmtsoc_litespimmap_bus_adr;
wire [31:0] mgmtsoc_litespimmap_bus_dat_w;
reg [31:0] mgmtsoc_litespimmap_bus_dat_r = 32'd0;
wire [3:0] mgmtsoc_litespimmap_bus_sel;
wire mgmtsoc_litespimmap_bus_cyc;
wire mgmtsoc_litespimmap_bus_stb;
reg mgmtsoc_litespimmap_bus_ack = 1'd0;
wire mgmtsoc_litespimmap_bus_we;
wire [2:0] mgmtsoc_litespimmap_bus_cti;
wire [1:0] mgmtsoc_litespimmap_bus_bte;
reg mgmtsoc_litespimmap_bus_err = 1'd0;
reg mgmtsoc_litespimmap_cs = 1'd0;
reg mgmtsoc_litespimmap_burst_cs = 1'd0;
reg [29:0] mgmtsoc_litespimmap_burst_adr = 30'd0;
reg mgmtsoc_litespimmap_wait = 1'd0;
wire mgmtsoc_litespimmap_done;
reg [8:0] mgmtsoc_litespimmap_count = 9'd256;
reg [7:0] mgmtsoc_litespimmap_storage = 8'd0;
reg mgmtsoc_litespimmap_re = 1'd0;
wire [7:0] mgmtsoc_litespimmap_spi_dummy_bits;
reg [31:0] mgmtsoc_litespimmap_dummy = 32'd57005;
reg [1:0] mgmtsoc_litespimmap = 2'd0;
wire mgmtsoc_port_mmap_user_port_source_valid;
wire mgmtsoc_port_mmap_user_port_source_ready;
wire mgmtsoc_port_mmap_user_port_source_first;
wire mgmtsoc_port_mmap_user_port_source_last;
wire [31:0] mgmtsoc_port_mmap_user_port_source_payload_data;
wire mgmtsoc_port_mmap_user_port_sink_valid;
wire mgmtsoc_port_mmap_user_port_sink_ready;
wire mgmtsoc_port_mmap_user_port_sink_first;
wire mgmtsoc_port_mmap_user_port_sink_last;
wire [31:0] mgmtsoc_port_mmap_user_port_sink_payload_data;
wire [5:0] mgmtsoc_port_mmap_user_port_sink_payload_len;
wire [3:0] mgmtsoc_port_mmap_user_port_sink_payload_width;
wire [7:0] mgmtsoc_port_mmap_user_port_sink_payload_mask;
wire mgmtsoc_port_mmap_internal_port_source_valid;
wire mgmtsoc_port_mmap_internal_port_source_ready;
wire mgmtsoc_port_mmap_internal_port_source_first;
wire mgmtsoc_port_mmap_internal_port_source_last;
wire [31:0] mgmtsoc_port_mmap_internal_port_source_payload_data;
wire mgmtsoc_port_mmap_internal_port_sink_valid;
wire mgmtsoc_port_mmap_internal_port_sink_ready;
wire mgmtsoc_port_mmap_internal_port_sink_first;
wire mgmtsoc_port_mmap_internal_port_sink_last;
wire [31:0] mgmtsoc_port_mmap_internal_port_sink_payload_data;
wire [5:0] mgmtsoc_port_mmap_internal_port_sink_payload_len;
wire [3:0] mgmtsoc_port_mmap_internal_port_sink_payload_width;
wire [7:0] mgmtsoc_port_mmap_internal_port_sink_payload_mask;
wire mgmtsoc_port_mmap_request;
wire mgmtsoc_master_sink_sink_valid;
wire mgmtsoc_master_sink_sink_ready;
wire mgmtsoc_master_sink_sink_first;
wire mgmtsoc_master_sink_sink_last;
wire [31:0] mgmtsoc_master_sink_sink_payload_data;
wire mgmtsoc_master_source_source_valid;
wire mgmtsoc_master_source_source_ready;
wire mgmtsoc_master_source_source_first;
wire mgmtsoc_master_source_source_last;
wire [31:0] mgmtsoc_master_source_source_payload_data;
wire [5:0] mgmtsoc_master_source_source_payload_len;
wire [3:0] mgmtsoc_master_source_source_payload_width;
wire [7:0] mgmtsoc_master_source_source_payload_mask;
wire mgmtsoc_master_cs;
reg mgmtsoc_master_cs_storage = 1'd0;
reg mgmtsoc_master_cs_re = 1'd0;
wire [7:0] mgmtsoc_master_len;
wire [3:0] mgmtsoc_master_width;
wire [7:0] mgmtsoc_master_mask;
reg [23:0] mgmtsoc_master_phyconfig_storage = 24'd0;
reg mgmtsoc_master_phyconfig_re = 1'd0;
reg mgmtsoc_master_rxtx_re = 1'd0;
wire [31:0] mgmtsoc_master_rxtx_r;
reg mgmtsoc_master_rxtx_we = 1'd0;
wire [31:0] mgmtsoc_master_rxtx_w;
wire mgmtsoc_master_tx_ready;
wire mgmtsoc_master_rx_ready;
reg [1:0] mgmtsoc_master_status_status = 2'd0;
wire mgmtsoc_master_status_we;
reg mgmtsoc_master_status_re = 1'd0;
wire mgmtsoc_master_tx_fifo_sink_valid;
wire mgmtsoc_master_tx_fifo_sink_ready;
reg mgmtsoc_master_tx_fifo_sink_first = 1'd0;
wire mgmtsoc_master_tx_fifo_sink_last;
wire [31:0] mgmtsoc_master_tx_fifo_sink_payload_data;
wire [5:0] mgmtsoc_master_tx_fifo_sink_payload_len;
wire [3:0] mgmtsoc_master_tx_fifo_sink_payload_width;
wire [7:0] mgmtsoc_master_tx_fifo_sink_payload_mask;
reg mgmtsoc_master_tx_fifo_source_valid = 1'd0;
wire mgmtsoc_master_tx_fifo_source_ready;
reg mgmtsoc_master_tx_fifo_source_first = 1'd0;
reg mgmtsoc_master_tx_fifo_source_last = 1'd0;
reg [31:0] mgmtsoc_master_tx_fifo_source_payload_data = 32'd0;
reg [5:0] mgmtsoc_master_tx_fifo_source_payload_len = 6'd0;
reg [3:0] mgmtsoc_master_tx_fifo_source_payload_width = 4'd0;
reg [7:0] mgmtsoc_master_tx_fifo_source_payload_mask = 8'd0;
wire mgmtsoc_master_rx_fifo_sink_valid;
wire mgmtsoc_master_rx_fifo_sink_ready;
wire mgmtsoc_master_rx_fifo_sink_first;
wire mgmtsoc_master_rx_fifo_sink_last;
wire [31:0] mgmtsoc_master_rx_fifo_sink_payload_data;
reg mgmtsoc_master_rx_fifo_source_valid = 1'd0;
wire mgmtsoc_master_rx_fifo_source_ready;
reg mgmtsoc_master_rx_fifo_source_first = 1'd0;
reg mgmtsoc_master_rx_fifo_source_last = 1'd0;
reg [31:0] mgmtsoc_master_rx_fifo_source_payload_data = 32'd0;
wire mgmtsoc_port_master_user_port_source_valid;
wire mgmtsoc_port_master_user_port_source_ready;
wire mgmtsoc_port_master_user_port_source_first;
wire mgmtsoc_port_master_user_port_source_last;
wire [31:0] mgmtsoc_port_master_user_port_source_payload_data;
wire mgmtsoc_port_master_user_port_sink_valid;
wire mgmtsoc_port_master_user_port_sink_ready;
wire mgmtsoc_port_master_user_port_sink_first;
wire mgmtsoc_port_master_user_port_sink_last;
wire [31:0] mgmtsoc_port_master_user_port_sink_payload_data;
wire [5:0] mgmtsoc_port_master_user_port_sink_payload_len;
wire [3:0] mgmtsoc_port_master_user_port_sink_payload_width;
wire [7:0] mgmtsoc_port_master_user_port_sink_payload_mask;
wire mgmtsoc_port_master_internal_port_source_valid;
wire mgmtsoc_port_master_internal_port_source_ready;
wire mgmtsoc_port_master_internal_port_source_first;
wire mgmtsoc_port_master_internal_port_source_last;
wire [31:0] mgmtsoc_port_master_internal_port_source_payload_data;
wire mgmtsoc_port_master_internal_port_sink_valid;
wire mgmtsoc_port_master_internal_port_sink_ready;
wire mgmtsoc_port_master_internal_port_sink_first;
wire mgmtsoc_port_master_internal_port_sink_last;
wire [31:0] mgmtsoc_port_master_internal_port_sink_payload_data;
wire [5:0] mgmtsoc_port_master_internal_port_sink_payload_len;
wire [3:0] mgmtsoc_port_master_internal_port_sink_payload_width;
wire [7:0] mgmtsoc_port_master_internal_port_sink_payload_mask;
wire mgmtsoc_port_master_request;
wire spi_master_start0;
wire [7:0] spi_master_length0;
reg spi_master_done0 = 1'd0;
reg spi_master_irq = 1'd0;
wire [7:0] spi_master_mosi;
reg [7:0] spi_master_miso = 8'd0;
wire spi_master_cs;
wire spi_master_cs_mode;
wire spi_master_loopback;
wire [15:0] spi_master_clk_divider0;
reg spi_master_start1 = 1'd0;
wire [7:0] spi_master_length1;
reg [15:0] spi_master_control_storage = 16'd0;
reg spi_master_control_re = 1'd0;
wire spi_master_done1;
wire spi_master_status_status;
wire spi_master_status_we;
reg spi_master_status_re = 1'd0;
reg [7:0] spi_master_mosi_storage = 8'd0;
reg spi_master_mosi_re = 1'd0;
wire [7:0] spi_master_miso_status;
wire spi_master_miso_we;
reg spi_master_miso_re = 1'd0;
wire spi_master_sel;
wire spi_master_mode0;
reg [16:0] spi_master_cs_storage = 17'd1;
reg spi_master_cs_re = 1'd0;
wire spi_master_mode1;
reg spi_master_loopback_storage = 1'd0;
reg spi_master_loopback_re = 1'd0;
reg spi_master_clk_enable = 1'd0;
reg spi_master_xfer_enable = 1'd0;
reg [2:0] spi_master_count = 3'd0;
reg spi_master_mosi_latch = 1'd0;
reg spi_master_miso_latch = 1'd0;
reg [15:0] spi_master_clk_divider1 = 16'd0;
wire spi_master_clk_rise;
wire spi_master_clk_fall;
reg [7:0] spi_master_mosi_data = 8'd0;
reg [2:0] spi_master_mosi_sel = 3'd0;
reg [7:0] spi_master_miso_data = 8'd0;
reg [15:0] spimaster_storage = 16'd100;
reg spimaster_re = 1'd0;
wire [29:0] mprj_adr;
wire [31:0] mprj_dat_w;
wire [31:0] mprj_dat_r;
wire [3:0] mprj_sel;
wire mprj_cyc;
wire mprj_stb;
wire mprj_ack;
wire mprj_we;
wire [2:0] mprj_cti;
wire [1:0] mprj_bte;
reg mprj_err = 1'd0;
reg mprj_wb_iena_storage = 1'd0;
reg mprj_wb_iena_re = 1'd0;
wire [29:0] hk_adr;
wire [31:0] hk_dat_w;
wire [31:0] hk_dat_r;
wire [3:0] hk_sel;
wire hk_cyc;
wire hk_stb;
wire hk_ack;
wire hk_we;
wire [2:0] hk_cti;
wire [1:0] hk_bte;
reg hk_err = 1'd0;
reg sys_uart_rx = 1'd0;
reg sys_uart_tx = 1'd1;
wire uart_phy_tx_sink_valid;
reg uart_phy_tx_sink_ready = 1'd0;
wire uart_phy_tx_sink_first;
wire uart_phy_tx_sink_last;
wire [7:0] uart_phy_tx_sink_payload_data;
reg [7:0] uart_phy_tx_data = 8'd0;
reg [3:0] uart_phy_tx_count = 4'd0;
reg uart_phy_tx_enable = 1'd0;
reg uart_phy_tx_tick = 1'd0;
reg [31:0] uart_phy_tx_phase = 32'd0;
reg uart_phy_rx_source_valid = 1'd0;
wire uart_phy_rx_source_ready;
reg uart_phy_rx_source_first = 1'd0;
reg uart_phy_rx_source_last = 1'd0;
reg [7:0] uart_phy_rx_source_payload_data = 8'd0;
reg [7:0] uart_phy_rx_data = 8'd0;
reg [3:0] uart_phy_rx_count = 4'd0;
reg uart_phy_rx_enable = 1'd0;
reg uart_phy_rx_tick = 1'd0;
reg [31:0] uart_phy_rx_phase = 32'd0;
wire uart_phy_rx_rx;
reg uart_phy_rx_rx_d = 1'd0;
reg uart_rxtx_re = 1'd0;
wire [7:0] uart_rxtx_r;
reg uart_rxtx_we = 1'd0;
wire [7:0] uart_rxtx_w;
wire uart_txfull_status;
wire uart_txfull_we;
reg uart_txfull_re = 1'd0;
wire uart_rxempty_status;
wire uart_rxempty_we;
reg uart_rxempty_re = 1'd0;
wire uart_irq;
wire uart_tx_status;
reg uart_tx_pending = 1'd0;
wire uart_tx_trigger;
reg uart_tx_clear = 1'd0;
reg uart_tx_trigger_d = 1'd0;
wire uart_rx_status;
reg uart_rx_pending = 1'd0;
wire uart_rx_trigger;
reg uart_rx_clear = 1'd0;
reg uart_rx_trigger_d = 1'd0;
wire uart_tx0;
wire uart_rx0;
reg [1:0] uart_status_status = 2'd0;
wire uart_status_we;
reg uart_status_re = 1'd0;
wire uart_tx1;
wire uart_rx1;
reg [1:0] uart_pending_status = 2'd0;
wire uart_pending_we;
reg uart_pending_re = 1'd0;
reg [1:0] uart_pending_r = 2'd0;
wire uart_tx2;
wire uart_rx2;
reg [1:0] uart_enable_storage = 2'd0;
reg uart_enable_re = 1'd0;
wire uart_txempty_status;
wire uart_txempty_we;
reg uart_txempty_re = 1'd0;
wire uart_rxfull_status;
wire uart_rxfull_we;
reg uart_rxfull_re = 1'd0;
wire uart_uart_sink_valid;
wire uart_uart_sink_ready;
wire uart_uart_sink_first;
wire uart_uart_sink_last;
wire [7:0] uart_uart_sink_payload_data;
wire uart_uart_source_valid;
wire uart_uart_source_ready;
wire uart_uart_source_first;
wire uart_uart_source_last;
wire [7:0] uart_uart_source_payload_data;
wire uart_tx_fifo_sink_valid;
wire uart_tx_fifo_sink_ready;
reg uart_tx_fifo_sink_first = 1'd0;
reg uart_tx_fifo_sink_last = 1'd0;
wire [7:0] uart_tx_fifo_sink_payload_data;
wire uart_tx_fifo_source_valid;
wire uart_tx_fifo_source_ready;
wire uart_tx_fifo_source_first;
wire uart_tx_fifo_source_last;
wire [7:0] uart_tx_fifo_source_payload_data;
wire uart_tx_fifo_re;
reg uart_tx_fifo_readable = 1'd0;
wire uart_tx_fifo_syncfifo_we;
wire uart_tx_fifo_syncfifo_writable;
wire uart_tx_fifo_syncfifo_re;
wire uart_tx_fifo_syncfifo_readable;
wire [9:0] uart_tx_fifo_syncfifo_din;
wire [9:0] uart_tx_fifo_syncfifo_dout;
reg [4:0] uart_tx_fifo_level0 = 5'd0;
reg uart_tx_fifo_replace = 1'd0;
reg [3:0] uart_tx_fifo_produce = 4'd0;
reg [3:0] uart_tx_fifo_consume = 4'd0;
reg [3:0] uart_tx_fifo_wrport_adr = 4'd0;
wire [9:0] uart_tx_fifo_wrport_dat_r;
wire uart_tx_fifo_wrport_we;
wire [9:0] uart_tx_fifo_wrport_dat_w;
wire uart_tx_fifo_do_read;
wire [3:0] uart_tx_fifo_rdport_adr;
wire [9:0] uart_tx_fifo_rdport_dat_r;
wire uart_tx_fifo_rdport_re;
wire [4:0] uart_tx_fifo_level1;
wire [7:0] uart_tx_fifo_fifo_in_payload_data;
wire uart_tx_fifo_fifo_in_first;
wire uart_tx_fifo_fifo_in_last;
wire [7:0] uart_tx_fifo_fifo_out_payload_data;
wire uart_tx_fifo_fifo_out_first;
wire uart_tx_fifo_fifo_out_last;
wire uart_rx_fifo_sink_valid;
wire uart_rx_fifo_sink_ready;
wire uart_rx_fifo_sink_first;
wire uart_rx_fifo_sink_last;
wire [7:0] uart_rx_fifo_sink_payload_data;
wire uart_rx_fifo_source_valid;
wire uart_rx_fifo_source_ready;
wire uart_rx_fifo_source_first;
wire uart_rx_fifo_source_last;
wire [7:0] uart_rx_fifo_source_payload_data;
wire uart_rx_fifo_re;
reg uart_rx_fifo_readable = 1'd0;
wire uart_rx_fifo_syncfifo_we;
wire uart_rx_fifo_syncfifo_writable;
wire uart_rx_fifo_syncfifo_re;
wire uart_rx_fifo_syncfifo_readable;
wire [9:0] uart_rx_fifo_syncfifo_din;
wire [9:0] uart_rx_fifo_syncfifo_dout;
reg [4:0] uart_rx_fifo_level0 = 5'd0;
reg uart_rx_fifo_replace = 1'd0;
reg [3:0] uart_rx_fifo_produce = 4'd0;
reg [3:0] uart_rx_fifo_consume = 4'd0;
reg [3:0] uart_rx_fifo_wrport_adr = 4'd0;
wire [9:0] uart_rx_fifo_wrport_dat_r;
wire uart_rx_fifo_wrport_we;
wire [9:0] uart_rx_fifo_wrport_dat_w;
wire uart_rx_fifo_do_read;
wire [3:0] uart_rx_fifo_rdport_adr;
wire [9:0] uart_rx_fifo_rdport_dat_r;
wire uart_rx_fifo_rdport_re;
wire [4:0] uart_rx_fifo_level1;
wire [7:0] uart_rx_fifo_fifo_in_payload_data;
wire uart_rx_fifo_fifo_in_first;
wire uart_rx_fifo_fifo_in_last;
wire [7:0] uart_rx_fifo_fifo_out_payload_data;
wire uart_rx_fifo_fifo_out_first;
wire uart_rx_fifo_fifo_out_last;
reg dbg_uart_dbg_uart_rx = 1'd0;
reg dbg_uart_dbg_uart_tx = 1'd1;
reg dbg_uart_tx_sink_valid = 1'd0;
reg dbg_uart_tx_sink_ready = 1'd0;
wire dbg_uart_tx_sink_last;
reg [7:0] dbg_uart_tx_sink_payload_data = 8'd0;
reg [7:0] dbg_uart_tx_data = 8'd0;
reg [3:0] dbg_uart_tx_count = 4'd0;
reg dbg_uart_tx_enable = 1'd0;
reg dbg_uart_tx_tick = 1'd0;
reg [31:0] dbg_uart_tx_phase = 32'd0;
reg dbg_uart_rx_source_valid = 1'd0;
reg dbg_uart_rx_source_ready = 1'd0;
reg [7:0] dbg_uart_rx_source_payload_data = 8'd0;
reg [7:0] dbg_uart_rx_data = 8'd0;
reg [3:0] dbg_uart_rx_count = 4'd0;
reg dbg_uart_rx_enable = 1'd0;
reg dbg_uart_rx_tick = 1'd0;
reg [31:0] dbg_uart_rx_phase = 32'd0;
wire dbg_uart_rx_rx;
reg dbg_uart_rx_rx_d = 1'd0;
wire [29:0] dbg_uart_wishbone_adr;
wire [31:0] dbg_uart_wishbone_dat_w;
wire [31:0] dbg_uart_wishbone_dat_r;
wire [3:0] dbg_uart_wishbone_sel;
reg dbg_uart_wishbone_cyc = 1'd0;
reg dbg_uart_wishbone_stb = 1'd0;
wire dbg_uart_wishbone_ack;
reg dbg_uart_wishbone_we = 1'd0;
reg [2:0] dbg_uart_wishbone_cti = 3'd0;
reg [1:0] dbg_uart_wishbone_bte = 2'd0;
wire dbg_uart_wishbone_err;
reg [7:0] dbg_uart_cmd = 8'd0;
reg dbg_uart_incr = 1'd0;
reg [7:0] dbg_uart_length = 8'd0;
reg [31:0] dbg_uart_address = 32'd0;
reg [31:0] dbg_uart_data = 32'd0;
reg [1:0] dbg_uart_bytes_count = 2'd0;
reg [7:0] dbg_uart_words_count = 8'd0;
wire dbg_uart_reset;
wire dbg_uart_wait;
wire dbg_uart_done;
reg [19:0] dbg_uart_count = 20'd1000000;
reg dbg_uart_is_ongoing = 1'd0;
reg debug_oeb_storage = 1'd0;
reg debug_oeb_re = 1'd0;
reg debug_mode_storage = 1'd0;
reg debug_mode_re = 1'd0;
wire uart_enabled_o;
reg uart_enabled_storage = 1'd0;
reg uart_enabled_re = 1'd0;
reg gpio_mode1_storage = 1'd0;
reg gpio_mode1_re = 1'd0;
reg gpio_mode0_storage = 1'd0;
reg gpio_mode0_re = 1'd0;
reg gpio_ien_storage = 1'd0;
reg gpio_ien_re = 1'd0;
reg gpio_oe_storage = 1'd0;
reg gpio_oe_re = 1'd0;
wire gpio_in_status;
wire gpio_in_we;
reg gpio_in_re = 1'd0;
reg gpio_out_storage = 1'd0;
reg gpio_out_re = 1'd0;
reg [127:0] la_ien_storage = 128'd0;
reg la_ien_re = 1'd0;
reg [127:0] la_oe_storage = 128'd0;
reg la_oe_re = 1'd0;
reg [127:0] la_in_status = 128'd0;
wire la_in_we;
reg la_in_re = 1'd0;
reg [127:0] la_out_storage = 128'd0;
reg la_out_re = 1'd0;
reg spi_enabled_storage = 1'd0;
reg spi_enabled_re = 1'd0;
reg [2:0] user_irq_ena_storage = 3'd0;
reg user_irq_ena_re = 1'd0;
wire gpioin0_in_status;
wire gpioin0_in_we;
reg gpioin0_in_re = 1'd0;
reg gpioin0_gpioin0_mode_storage = 1'd0;
reg gpioin0_gpioin0_mode_re = 1'd0;
reg gpioin0_gpioin0_edge_storage = 1'd0;
reg gpioin0_gpioin0_edge_re = 1'd0;
wire gpioin0_gpioin0_irq;
reg gpioin0_gpioin0_in_pads_n_d = 1'd0;
wire gpioin0_gpioin0_status;
reg gpioin0_gpioin0_pending = 1'd0;
reg gpioin0_gpioin0_trigger = 1'd0;
reg gpioin0_gpioin0_clear = 1'd0;
reg gpioin0_gpioin0_trigger_d = 1'd0;
wire gpioin1_in_status;
wire gpioin1_in_we;
reg gpioin1_in_re = 1'd0;
reg gpioin1_gpioin1_mode_storage = 1'd0;
reg gpioin1_gpioin1_mode_re = 1'd0;
reg gpioin1_gpioin1_edge_storage = 1'd0;
reg gpioin1_gpioin1_edge_re = 1'd0;
wire gpioin1_gpioin1_irq;
reg gpioin1_gpioin1_in_pads_n_d = 1'd0;
wire gpioin1_gpioin1_status;
reg gpioin1_gpioin1_pending = 1'd0;
reg gpioin1_gpioin1_trigger = 1'd0;
reg gpioin1_gpioin1_clear = 1'd0;
reg gpioin1_gpioin1_trigger_d = 1'd0;
wire gpioin2_in_status;
wire gpioin2_in_we;
reg gpioin2_in_re = 1'd0;
reg gpioin2_gpioin2_mode_storage = 1'd0;
reg gpioin2_gpioin2_mode_re = 1'd0;
reg gpioin2_gpioin2_edge_storage = 1'd0;
reg gpioin2_gpioin2_edge_re = 1'd0;
wire gpioin2_gpioin2_irq;
reg gpioin2_gpioin2_in_pads_n_d = 1'd0;
wire gpioin2_gpioin2_status;
reg gpioin2_gpioin2_pending = 1'd0;
reg gpioin2_gpioin2_trigger = 1'd0;
reg gpioin2_gpioin2_clear = 1'd0;
reg gpioin2_gpioin2_trigger_d = 1'd0;
wire gpioin3_in_status;
wire gpioin3_in_we;
reg gpioin3_in_re = 1'd0;
reg gpioin3_gpioin3_mode_storage = 1'd0;
reg gpioin3_gpioin3_mode_re = 1'd0;
reg gpioin3_gpioin3_edge_storage = 1'd0;
reg gpioin3_gpioin3_edge_re = 1'd0;
wire gpioin3_gpioin3_irq;
reg gpioin3_gpioin3_in_pads_n_d = 1'd0;
wire gpioin3_gpioin3_status;
reg gpioin3_gpioin3_pending = 1'd0;
reg gpioin3_gpioin3_trigger = 1'd0;
reg gpioin3_gpioin3_clear = 1'd0;
reg gpioin3_gpioin3_trigger_d = 1'd0;
wire gpioin4_in_status;
wire gpioin4_in_we;
reg gpioin4_in_re = 1'd0;
reg gpioin4_gpioin4_mode_storage = 1'd0;
reg gpioin4_gpioin4_mode_re = 1'd0;
reg gpioin4_gpioin4_edge_storage = 1'd0;
reg gpioin4_gpioin4_edge_re = 1'd0;
wire gpioin4_gpioin4_irq;
reg gpioin4_gpioin4_in_pads_n_d = 1'd0;
wire gpioin4_gpioin4_status;
reg gpioin4_gpioin4_pending = 1'd0;
reg gpioin4_gpioin4_trigger = 1'd0;
reg gpioin4_gpioin4_clear = 1'd0;
reg gpioin4_gpioin4_trigger_d = 1'd0;
wire gpioin5_in_status;
wire gpioin5_in_we;
reg gpioin5_in_re = 1'd0;
reg gpioin5_gpioin5_mode_storage = 1'd0;
reg gpioin5_gpioin5_mode_re = 1'd0;
reg gpioin5_gpioin5_edge_storage = 1'd0;
reg gpioin5_gpioin5_edge_re = 1'd0;
wire gpioin5_gpioin5_irq;
reg gpioin5_gpioin5_in_pads_n_d = 1'd0;
wire gpioin5_gpioin5_status;
reg gpioin5_gpioin5_pending = 1'd0;
reg gpioin5_gpioin5_trigger = 1'd0;
reg gpioin5_gpioin5_clear = 1'd0;
reg gpioin5_gpioin5_trigger_d = 1'd0;
reg [1:0] litespiphy_state = 2'd0;
reg [1:0] litespiphy_next_state = 2'd0;
reg [7:0] mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value = 8'd0;
reg mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce = 1'd0;
wire [1:0] litespi_request;
reg litespi_grant = 1'd0;
reg litespi_tx_mux_source_valid = 1'd0;
wire litespi_tx_mux_source_ready;
reg litespi_tx_mux_source_first = 1'd0;
reg litespi_tx_mux_source_last = 1'd0;
reg [31:0] litespi_tx_mux_source_payload_data = 32'd0;
reg [5:0] litespi_tx_mux_source_payload_len = 6'd0;
reg [3:0] litespi_tx_mux_source_payload_width = 4'd0;
reg [7:0] litespi_tx_mux_source_payload_mask = 8'd0;
wire litespi_tx_mux_endpoint0_sink_valid;
reg litespi_tx_mux_endpoint0_sink_ready = 1'd0;
wire litespi_tx_mux_endpoint0_sink_first;
wire litespi_tx_mux_endpoint0_sink_last;
wire [31:0] litespi_tx_mux_endpoint0_sink_payload_data;
wire [5:0] litespi_tx_mux_endpoint0_sink_payload_len;
wire [3:0] litespi_tx_mux_endpoint0_sink_payload_width;
wire [7:0] litespi_tx_mux_endpoint0_sink_payload_mask;
wire litespi_tx_mux_endpoint1_sink_valid;
reg litespi_tx_mux_endpoint1_sink_ready = 1'd0;
wire litespi_tx_mux_endpoint1_sink_first;
wire litespi_tx_mux_endpoint1_sink_last;
wire [31:0] litespi_tx_mux_endpoint1_sink_payload_data;
wire [5:0] litespi_tx_mux_endpoint1_sink_payload_len;
wire [3:0] litespi_tx_mux_endpoint1_sink_payload_width;
wire [7:0] litespi_tx_mux_endpoint1_sink_payload_mask;
wire litespi_tx_mux_sel;
wire litespi_rx_demux_sink_valid;
reg litespi_rx_demux_sink_ready = 1'd0;
wire litespi_rx_demux_sink_first;
wire litespi_rx_demux_sink_last;
wire [31:0] litespi_rx_demux_sink_payload_data;
reg litespi_rx_demux_endpoint0_source_valid = 1'd0;
wire litespi_rx_demux_endpoint0_source_ready;
reg litespi_rx_demux_endpoint0_source_first = 1'd0;
reg litespi_rx_demux_endpoint0_source_last = 1'd0;
reg [31:0] litespi_rx_demux_endpoint0_source_payload_data = 32'd0;
reg litespi_rx_demux_endpoint1_source_valid = 1'd0;
wire litespi_rx_demux_endpoint1_source_ready;
reg litespi_rx_demux_endpoint1_source_first = 1'd0;
reg litespi_rx_demux_endpoint1_source_last = 1'd0;
reg [31:0] litespi_rx_demux_endpoint1_source_payload_data = 32'd0;
wire litespi_rx_demux_sel;
reg [3:0] litespi_state = 4'd0;
reg [3:0] litespi_next_state = 4'd0;
reg mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = 1'd0;
reg mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd0;
reg [29:0] mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = 30'd0;
reg mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd0;
reg [1:0] spimaster_state = 2'd0;
reg [1:0] spimaster_next_state = 2'd0;
reg [2:0] spi_master_count_spimaster_next_value = 3'd0;
reg spi_master_count_spimaster_next_value_ce = 1'd0;
reg rs232phy_rs232phytx_state = 1'd0;
reg rs232phy_rs232phytx_next_state = 1'd0;
reg [3:0] uart_phy_tx_count_rs232phy_rs232phytx_next_value0 = 4'd0;
reg uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0 = 1'd0;
reg sys_uart_tx_rs232phy_rs232phytx_next_value1 = 1'd0;
reg sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd0;
reg [7:0] uart_phy_tx_data_rs232phy_rs232phytx_next_value2 = 8'd0;
reg uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2 = 1'd0;
reg rs232phy_rs232phyrx_state = 1'd0;
reg rs232phy_rs232phyrx_next_state = 1'd0;
reg [3:0] uart_phy_rx_count_rs232phy_rs232phyrx_next_value0 = 4'd0;
reg uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0 = 1'd0;
reg [7:0] uart_phy_rx_data_rs232phy_rs232phyrx_next_value1 = 8'd0;
reg uart_phy_rx_data_rs232phy_rs232phyrx_next_value_ce1 = 1'd0;
reg uartwishbonebridge_rs232phytx_state = 1'd0;
reg uartwishbonebridge_rs232phytx_next_state = 1'd0;
reg [3:0] dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0 = 4'd0;
reg dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0 = 1'd0;
reg dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = 1'd0;
reg dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd0;
reg [7:0] dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2 = 8'd0;
reg dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2 = 1'd0;
reg uartwishbonebridge_rs232phyrx_state = 1'd0;
reg uartwishbonebridge_rs232phyrx_next_state = 1'd0;
reg [3:0] dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0 = 4'd0;
reg dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0 = 1'd0;
reg [7:0] dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value1 = 8'd0;
reg dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value_ce1 = 1'd0;
reg [2:0] uartwishbonebridge_state = 3'd0;
reg [2:0] uartwishbonebridge_next_state = 3'd0;
reg [1:0] dbg_uart_bytes_count_uartwishbonebridge_next_value0 = 2'd0;
reg dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd0;
reg [7:0] dbg_uart_words_count_uartwishbonebridge_next_value1 = 8'd0;
reg dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd0;
reg [7:0] dbg_uart_cmd_uartwishbonebridge_next_value2 = 8'd0;
reg dbg_uart_cmd_uartwishbonebridge_next_value_ce2 = 1'd0;
reg [7:0] dbg_uart_length_uartwishbonebridge_next_value3 = 8'd0;
reg dbg_uart_length_uartwishbonebridge_next_value_ce3 = 1'd0;
reg [31:0] dbg_uart_address_uartwishbonebridge_next_value4 = 32'd0;
reg dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd0;
reg dbg_uart_incr_uartwishbonebridge_next_value5 = 1'd0;
reg dbg_uart_incr_uartwishbonebridge_next_value_ce5 = 1'd0;
reg [31:0] dbg_uart_data_uartwishbonebridge_next_value6 = 32'd0;
reg dbg_uart_data_uartwishbonebridge_next_value_ce6 = 1'd0;
wire gpioin0_i00;
wire gpioin0_status_status;
wire gpioin0_status_we;
reg gpioin0_status_re = 1'd0;
wire gpioin0_i01;
wire gpioin0_pending_status;
wire gpioin0_pending_we;
reg gpioin0_pending_re = 1'd0;
reg gpioin0_pending_r = 1'd0;
wire gpioin0_i02;
reg gpioin0_enable_storage = 1'd0;
reg gpioin0_enable_re = 1'd0;
wire gpioin1_i00;
wire gpioin1_status_status;
wire gpioin1_status_we;
reg gpioin1_status_re = 1'd0;
wire gpioin1_i01;
wire gpioin1_pending_status;
wire gpioin1_pending_we;
reg gpioin1_pending_re = 1'd0;
reg gpioin1_pending_r = 1'd0;
wire gpioin1_i02;
reg gpioin1_enable_storage = 1'd0;
reg gpioin1_enable_re = 1'd0;
wire gpioin2_i00;
wire gpioin2_status_status;
wire gpioin2_status_we;
reg gpioin2_status_re = 1'd0;
wire gpioin2_i01;
wire gpioin2_pending_status;
wire gpioin2_pending_we;
reg gpioin2_pending_re = 1'd0;
reg gpioin2_pending_r = 1'd0;
wire gpioin2_i02;
reg gpioin2_enable_storage = 1'd0;
reg gpioin2_enable_re = 1'd0;
wire gpioin3_i00;
wire gpioin3_status_status;
wire gpioin3_status_we;
reg gpioin3_status_re = 1'd0;
wire gpioin3_i01;
wire gpioin3_pending_status;
wire gpioin3_pending_we;
reg gpioin3_pending_re = 1'd0;
reg gpioin3_pending_r = 1'd0;
wire gpioin3_i02;
reg gpioin3_enable_storage = 1'd0;
reg gpioin3_enable_re = 1'd0;
wire gpioin4_i00;
wire gpioin4_status_status;
wire gpioin4_status_we;
reg gpioin4_status_re = 1'd0;
wire gpioin4_i01;
wire gpioin4_pending_status;
wire gpioin4_pending_we;
reg gpioin4_pending_re = 1'd0;
reg gpioin4_pending_r = 1'd0;
wire gpioin4_i02;
reg gpioin4_enable_storage = 1'd0;
reg gpioin4_enable_re = 1'd0;
wire gpioin5_i00;
wire gpioin5_status_status;
wire gpioin5_status_we;
reg gpioin5_status_re = 1'd0;
wire gpioin5_i01;
wire gpioin5_pending_status;
wire gpioin5_pending_we;
reg gpioin5_pending_re = 1'd0;
reg gpioin5_pending_r = 1'd0;
wire gpioin5_i02;
reg gpioin5_enable_storage = 1'd0;
reg gpioin5_enable_re = 1'd0;
reg [13:0] mgmtsoc_adr = 14'd0;
reg mgmtsoc_we = 1'd0;
reg [31:0] mgmtsoc_dat_w = 32'd0;
wire [31:0] mgmtsoc_dat_r;
wire [29:0] mgmtsoc_wishbone_adr;
wire [31:0] mgmtsoc_wishbone_dat_w;
reg [31:0] mgmtsoc_wishbone_dat_r = 32'd0;
wire [3:0] mgmtsoc_wishbone_sel;
wire mgmtsoc_wishbone_cyc;
wire mgmtsoc_wishbone_stb;
reg mgmtsoc_wishbone_ack = 1'd0;
wire mgmtsoc_wishbone_we;
wire [2:0] mgmtsoc_wishbone_cti;
wire [1:0] mgmtsoc_wishbone_bte;
reg mgmtsoc_wishbone_err = 1'd0;
wire [29:0] shared_adr;
wire [31:0] shared_dat_w;
reg [31:0] shared_dat_r = 32'd0;
wire [3:0] shared_sel;
wire shared_cyc;
wire shared_stb;
reg shared_ack = 1'd0;
wire shared_we;
wire [2:0] shared_cti;
wire [1:0] shared_bte;
wire shared_err;
wire [2:0] request;
reg [1:0] grant = 2'd0;
reg [6:0] slave_sel = 7'd0;
reg [6:0] slave_sel_r = 7'd0;
reg error = 1'd0;
wire wait_1;
wire done;
reg [19:0] count = 20'd1000000;
wire [13:0] interface0_bank_bus_adr;
wire interface0_bank_bus_we;
wire [31:0] interface0_bank_bus_dat_w;
reg [31:0] interface0_bank_bus_dat_r = 32'd0;
reg csrbank0_reset0_re = 1'd0;
wire [1:0] csrbank0_reset0_r;
reg csrbank0_reset0_we = 1'd0;
wire [1:0] csrbank0_reset0_w;
reg csrbank0_scratch0_re = 1'd0;
wire [31:0] csrbank0_scratch0_r;
reg csrbank0_scratch0_we = 1'd0;
wire [31:0] csrbank0_scratch0_w;
reg csrbank0_bus_errors_re = 1'd0;
wire [31:0] csrbank0_bus_errors_r;
reg csrbank0_bus_errors_we = 1'd0;
wire [31:0] csrbank0_bus_errors_w;
wire csrbank0_sel;
wire [13:0] interface1_bank_bus_adr;
wire interface1_bank_bus_we;
wire [31:0] interface1_bank_bus_dat_w;
reg [31:0] interface1_bank_bus_dat_r = 32'd0;
reg csrbank1_out0_re = 1'd0;
wire csrbank1_out0_r;
reg csrbank1_out0_we = 1'd0;
wire csrbank1_out0_w;
wire csrbank1_sel;
wire [13:0] interface2_bank_bus_adr;
wire interface2_bank_bus_we;
wire [31:0] interface2_bank_bus_dat_w;
reg [31:0] interface2_bank_bus_dat_r = 32'd0;
reg csrbank2_out0_re = 1'd0;
wire csrbank2_out0_r;
reg csrbank2_out0_we = 1'd0;
wire csrbank2_out0_w;
wire csrbank2_sel;
wire [13:0] interface3_bank_bus_adr;
wire interface3_bank_bus_we;
wire [31:0] interface3_bank_bus_dat_w;
reg [31:0] interface3_bank_bus_dat_r = 32'd0;
reg csrbank3_mmap_dummy_bits0_re = 1'd0;
wire [7:0] csrbank3_mmap_dummy_bits0_r;
reg csrbank3_mmap_dummy_bits0_we = 1'd0;
wire [7:0] csrbank3_mmap_dummy_bits0_w;
reg csrbank3_master_cs0_re = 1'd0;
wire csrbank3_master_cs0_r;
reg csrbank3_master_cs0_we = 1'd0;
wire csrbank3_master_cs0_w;
reg csrbank3_master_phyconfig0_re = 1'd0;
wire [23:0] csrbank3_master_phyconfig0_r;
reg csrbank3_master_phyconfig0_we = 1'd0;
wire [23:0] csrbank3_master_phyconfig0_w;
reg csrbank3_master_status_re = 1'd0;
wire [1:0] csrbank3_master_status_r;
reg csrbank3_master_status_we = 1'd0;
wire [1:0] csrbank3_master_status_w;
wire csrbank3_sel;
wire [13:0] interface4_bank_bus_adr;
wire interface4_bank_bus_we;
wire [31:0] interface4_bank_bus_dat_w;
reg [31:0] interface4_bank_bus_dat_r = 32'd0;
reg csrbank4_clk_divisor0_re = 1'd0;
wire [7:0] csrbank4_clk_divisor0_r;
reg csrbank4_clk_divisor0_we = 1'd0;
wire [7:0] csrbank4_clk_divisor0_w;
wire csrbank4_sel;
wire [13:0] interface5_bank_bus_adr;
wire interface5_bank_bus_we;
wire [31:0] interface5_bank_bus_dat_w;
reg [31:0] interface5_bank_bus_dat_r = 32'd0;
reg csrbank5_mode10_re = 1'd0;
wire csrbank5_mode10_r;
reg csrbank5_mode10_we = 1'd0;
wire csrbank5_mode10_w;
reg csrbank5_mode00_re = 1'd0;
wire csrbank5_mode00_r;
reg csrbank5_mode00_we = 1'd0;
wire csrbank5_mode00_w;
reg csrbank5_ien0_re = 1'd0;
wire csrbank5_ien0_r;
reg csrbank5_ien0_we = 1'd0;
wire csrbank5_ien0_w;
reg csrbank5_oe0_re = 1'd0;
wire csrbank5_oe0_r;
reg csrbank5_oe0_we = 1'd0;
wire csrbank5_oe0_w;
reg csrbank5_in_re = 1'd0;
wire csrbank5_in_r;
reg csrbank5_in_we = 1'd0;
wire csrbank5_in_w;
reg csrbank5_out0_re = 1'd0;
wire csrbank5_out0_r;
reg csrbank5_out0_we = 1'd0;
wire csrbank5_out0_w;
wire csrbank5_sel;
wire [13:0] interface6_bank_bus_adr;
wire interface6_bank_bus_we;
wire [31:0] interface6_bank_bus_dat_w;
reg [31:0] interface6_bank_bus_dat_r = 32'd0;
reg csrbank6_ien3_re = 1'd0;
wire [31:0] csrbank6_ien3_r;
reg csrbank6_ien3_we = 1'd0;
wire [31:0] csrbank6_ien3_w;
reg csrbank6_ien2_re = 1'd0;
wire [31:0] csrbank6_ien2_r;
reg csrbank6_ien2_we = 1'd0;
wire [31:0] csrbank6_ien2_w;
reg csrbank6_ien1_re = 1'd0;
wire [31:0] csrbank6_ien1_r;
reg csrbank6_ien1_we = 1'd0;
wire [31:0] csrbank6_ien1_w;
reg csrbank6_ien0_re = 1'd0;
wire [31:0] csrbank6_ien0_r;
reg csrbank6_ien0_we = 1'd0;
wire [31:0] csrbank6_ien0_w;
reg csrbank6_oe3_re = 1'd0;
wire [31:0] csrbank6_oe3_r;
reg csrbank6_oe3_we = 1'd0;
wire [31:0] csrbank6_oe3_w;
reg csrbank6_oe2_re = 1'd0;
wire [31:0] csrbank6_oe2_r;
reg csrbank6_oe2_we = 1'd0;
wire [31:0] csrbank6_oe2_w;
reg csrbank6_oe1_re = 1'd0;
wire [31:0] csrbank6_oe1_r;
reg csrbank6_oe1_we = 1'd0;
wire [31:0] csrbank6_oe1_w;
reg csrbank6_oe0_re = 1'd0;
wire [31:0] csrbank6_oe0_r;
reg csrbank6_oe0_we = 1'd0;
wire [31:0] csrbank6_oe0_w;
reg csrbank6_in3_re = 1'd0;
wire [31:0] csrbank6_in3_r;
reg csrbank6_in3_we = 1'd0;
wire [31:0] csrbank6_in3_w;
reg csrbank6_in2_re = 1'd0;
wire [31:0] csrbank6_in2_r;
reg csrbank6_in2_we = 1'd0;
wire [31:0] csrbank6_in2_w;
reg csrbank6_in1_re = 1'd0;
wire [31:0] csrbank6_in1_r;
reg csrbank6_in1_we = 1'd0;
wire [31:0] csrbank6_in1_w;
reg csrbank6_in0_re = 1'd0;
wire [31:0] csrbank6_in0_r;
reg csrbank6_in0_we = 1'd0;
wire [31:0] csrbank6_in0_w;
reg csrbank6_out3_re = 1'd0;
wire [31:0] csrbank6_out3_r;
reg csrbank6_out3_we = 1'd0;
wire [31:0] csrbank6_out3_w;
reg csrbank6_out2_re = 1'd0;
wire [31:0] csrbank6_out2_r;
reg csrbank6_out2_we = 1'd0;
wire [31:0] csrbank6_out2_w;
reg csrbank6_out1_re = 1'd0;
wire [31:0] csrbank6_out1_r;
reg csrbank6_out1_we = 1'd0;
wire [31:0] csrbank6_out1_w;
reg csrbank6_out0_re = 1'd0;
wire [31:0] csrbank6_out0_r;
reg csrbank6_out0_we = 1'd0;
wire [31:0] csrbank6_out0_w;
wire csrbank6_sel;
wire [13:0] interface7_bank_bus_adr;
wire interface7_bank_bus_we;
wire [31:0] interface7_bank_bus_dat_w;
reg [31:0] interface7_bank_bus_dat_r = 32'd0;
reg csrbank7_out0_re = 1'd0;
wire csrbank7_out0_r;
reg csrbank7_out0_we = 1'd0;
wire csrbank7_out0_w;
wire csrbank7_sel;
wire [13:0] interface8_bank_bus_adr;
wire interface8_bank_bus_we;
wire [31:0] interface8_bank_bus_dat_w;
reg [31:0] interface8_bank_bus_dat_r = 32'd0;
reg csrbank8_out0_re = 1'd0;
wire csrbank8_out0_r;
reg csrbank8_out0_we = 1'd0;
wire csrbank8_out0_w;
wire csrbank8_sel;
wire [13:0] interface9_bank_bus_adr;
wire interface9_bank_bus_we;
wire [31:0] interface9_bank_bus_dat_w;
reg [31:0] interface9_bank_bus_dat_r = 32'd0;
reg csrbank9_control0_re = 1'd0;
wire [15:0] csrbank9_control0_r;
reg csrbank9_control0_we = 1'd0;
wire [15:0] csrbank9_control0_w;
reg csrbank9_status_re = 1'd0;
wire csrbank9_status_r;
reg csrbank9_status_we = 1'd0;
wire csrbank9_status_w;
reg csrbank9_mosi0_re = 1'd0;
wire [7:0] csrbank9_mosi0_r;
reg csrbank9_mosi0_we = 1'd0;
wire [7:0] csrbank9_mosi0_w;
reg csrbank9_miso_re = 1'd0;
wire [7:0] csrbank9_miso_r;
reg csrbank9_miso_we = 1'd0;
wire [7:0] csrbank9_miso_w;
reg csrbank9_cs0_re = 1'd0;
wire [16:0] csrbank9_cs0_r;
reg csrbank9_cs0_we = 1'd0;
wire [16:0] csrbank9_cs0_w;
reg csrbank9_loopback0_re = 1'd0;
wire csrbank9_loopback0_r;
reg csrbank9_loopback0_we = 1'd0;
wire csrbank9_loopback0_w;
reg csrbank9_clk_divider0_re = 1'd0;
wire [15:0] csrbank9_clk_divider0_r;
reg csrbank9_clk_divider0_we = 1'd0;
wire [15:0] csrbank9_clk_divider0_w;
wire csrbank9_sel;
wire [13:0] interface10_bank_bus_adr;
wire interface10_bank_bus_we;
wire [31:0] interface10_bank_bus_dat_w;
reg [31:0] interface10_bank_bus_dat_r = 32'd0;
reg csrbank10_load0_re = 1'd0;
wire [31:0] csrbank10_load0_r;
reg csrbank10_load0_we = 1'd0;
wire [31:0] csrbank10_load0_w;
reg csrbank10_reload0_re = 1'd0;
wire [31:0] csrbank10_reload0_r;
reg csrbank10_reload0_we = 1'd0;
wire [31:0] csrbank10_reload0_w;
reg csrbank10_en0_re = 1'd0;
wire csrbank10_en0_r;
reg csrbank10_en0_we = 1'd0;
wire csrbank10_en0_w;
reg csrbank10_update_value0_re = 1'd0;
wire csrbank10_update_value0_r;
reg csrbank10_update_value0_we = 1'd0;
wire csrbank10_update_value0_w;
reg csrbank10_value_re = 1'd0;
wire [31:0] csrbank10_value_r;
reg csrbank10_value_we = 1'd0;
wire [31:0] csrbank10_value_w;
reg csrbank10_ev_status_re = 1'd0;
wire csrbank10_ev_status_r;
reg csrbank10_ev_status_we = 1'd0;
wire csrbank10_ev_status_w;
reg csrbank10_ev_pending_re = 1'd0;
wire csrbank10_ev_pending_r;
reg csrbank10_ev_pending_we = 1'd0;
wire csrbank10_ev_pending_w;
reg csrbank10_ev_enable0_re = 1'd0;
wire csrbank10_ev_enable0_r;
reg csrbank10_ev_enable0_we = 1'd0;
wire csrbank10_ev_enable0_w;
wire csrbank10_sel;
wire [13:0] interface11_bank_bus_adr;
wire interface11_bank_bus_we;
wire [31:0] interface11_bank_bus_dat_w;
reg [31:0] interface11_bank_bus_dat_r = 32'd0;
reg csrbank11_txfull_re = 1'd0;
wire csrbank11_txfull_r;
reg csrbank11_txfull_we = 1'd0;
wire csrbank11_txfull_w;
reg csrbank11_rxempty_re = 1'd0;
wire csrbank11_rxempty_r;
reg csrbank11_rxempty_we = 1'd0;
wire csrbank11_rxempty_w;
reg csrbank11_ev_status_re = 1'd0;
wire [1:0] csrbank11_ev_status_r;
reg csrbank11_ev_status_we = 1'd0;
wire [1:0] csrbank11_ev_status_w;
reg csrbank11_ev_pending_re = 1'd0;
wire [1:0] csrbank11_ev_pending_r;
reg csrbank11_ev_pending_we = 1'd0;
wire [1:0] csrbank11_ev_pending_w;
reg csrbank11_ev_enable0_re = 1'd0;
wire [1:0] csrbank11_ev_enable0_r;
reg csrbank11_ev_enable0_we = 1'd0;
wire [1:0] csrbank11_ev_enable0_w;
reg csrbank11_txempty_re = 1'd0;
wire csrbank11_txempty_r;
reg csrbank11_txempty_we = 1'd0;
wire csrbank11_txempty_w;
reg csrbank11_rxfull_re = 1'd0;
wire csrbank11_rxfull_r;
reg csrbank11_rxfull_we = 1'd0;
wire csrbank11_rxfull_w;
wire csrbank11_sel;
wire [13:0] interface12_bank_bus_adr;
wire interface12_bank_bus_we;
wire [31:0] interface12_bank_bus_dat_w;
reg [31:0] interface12_bank_bus_dat_r = 32'd0;
reg csrbank12_out0_re = 1'd0;
wire csrbank12_out0_r;
reg csrbank12_out0_we = 1'd0;
wire csrbank12_out0_w;
wire csrbank12_sel;
wire [13:0] interface13_bank_bus_adr;
wire interface13_bank_bus_we;
wire [31:0] interface13_bank_bus_dat_w;
reg [31:0] interface13_bank_bus_dat_r = 32'd0;
reg csrbank13_in_re = 1'd0;
wire csrbank13_in_r;
reg csrbank13_in_we = 1'd0;
wire csrbank13_in_w;
reg csrbank13_mode0_re = 1'd0;
wire csrbank13_mode0_r;
reg csrbank13_mode0_we = 1'd0;
wire csrbank13_mode0_w;
reg csrbank13_edge0_re = 1'd0;
wire csrbank13_edge0_r;
reg csrbank13_edge0_we = 1'd0;
wire csrbank13_edge0_w;
reg csrbank13_ev_status_re = 1'd0;
wire csrbank13_ev_status_r;
reg csrbank13_ev_status_we = 1'd0;
wire csrbank13_ev_status_w;
reg csrbank13_ev_pending_re = 1'd0;
wire csrbank13_ev_pending_r;
reg csrbank13_ev_pending_we = 1'd0;
wire csrbank13_ev_pending_w;
reg csrbank13_ev_enable0_re = 1'd0;
wire csrbank13_ev_enable0_r;
reg csrbank13_ev_enable0_we = 1'd0;
wire csrbank13_ev_enable0_w;
wire csrbank13_sel;
wire [13:0] interface14_bank_bus_adr;
wire interface14_bank_bus_we;
wire [31:0] interface14_bank_bus_dat_w;
reg [31:0] interface14_bank_bus_dat_r = 32'd0;
reg csrbank14_in_re = 1'd0;
wire csrbank14_in_r;
reg csrbank14_in_we = 1'd0;
wire csrbank14_in_w;
reg csrbank14_mode0_re = 1'd0;
wire csrbank14_mode0_r;
reg csrbank14_mode0_we = 1'd0;
wire csrbank14_mode0_w;
reg csrbank14_edge0_re = 1'd0;
wire csrbank14_edge0_r;
reg csrbank14_edge0_we = 1'd0;
wire csrbank14_edge0_w;
reg csrbank14_ev_status_re = 1'd0;
wire csrbank14_ev_status_r;
reg csrbank14_ev_status_we = 1'd0;
wire csrbank14_ev_status_w;
reg csrbank14_ev_pending_re = 1'd0;
wire csrbank14_ev_pending_r;
reg csrbank14_ev_pending_we = 1'd0;
wire csrbank14_ev_pending_w;
reg csrbank14_ev_enable0_re = 1'd0;
wire csrbank14_ev_enable0_r;
reg csrbank14_ev_enable0_we = 1'd0;
wire csrbank14_ev_enable0_w;
wire csrbank14_sel;
wire [13:0] interface15_bank_bus_adr;
wire interface15_bank_bus_we;
wire [31:0] interface15_bank_bus_dat_w;
reg [31:0] interface15_bank_bus_dat_r = 32'd0;
reg csrbank15_in_re = 1'd0;
wire csrbank15_in_r;
reg csrbank15_in_we = 1'd0;
wire csrbank15_in_w;
reg csrbank15_mode0_re = 1'd0;
wire csrbank15_mode0_r;
reg csrbank15_mode0_we = 1'd0;
wire csrbank15_mode0_w;
reg csrbank15_edge0_re = 1'd0;
wire csrbank15_edge0_r;
reg csrbank15_edge0_we = 1'd0;
wire csrbank15_edge0_w;
reg csrbank15_ev_status_re = 1'd0;
wire csrbank15_ev_status_r;
reg csrbank15_ev_status_we = 1'd0;
wire csrbank15_ev_status_w;
reg csrbank15_ev_pending_re = 1'd0;
wire csrbank15_ev_pending_r;
reg csrbank15_ev_pending_we = 1'd0;
wire csrbank15_ev_pending_w;
reg csrbank15_ev_enable0_re = 1'd0;
wire csrbank15_ev_enable0_r;
reg csrbank15_ev_enable0_we = 1'd0;
wire csrbank15_ev_enable0_w;
wire csrbank15_sel;
wire [13:0] interface16_bank_bus_adr;
wire interface16_bank_bus_we;
wire [31:0] interface16_bank_bus_dat_w;
reg [31:0] interface16_bank_bus_dat_r = 32'd0;
reg csrbank16_in_re = 1'd0;
wire csrbank16_in_r;
reg csrbank16_in_we = 1'd0;
wire csrbank16_in_w;
reg csrbank16_mode0_re = 1'd0;
wire csrbank16_mode0_r;
reg csrbank16_mode0_we = 1'd0;
wire csrbank16_mode0_w;
reg csrbank16_edge0_re = 1'd0;
wire csrbank16_edge0_r;
reg csrbank16_edge0_we = 1'd0;
wire csrbank16_edge0_w;
reg csrbank16_ev_status_re = 1'd0;
wire csrbank16_ev_status_r;
reg csrbank16_ev_status_we = 1'd0;
wire csrbank16_ev_status_w;
reg csrbank16_ev_pending_re = 1'd0;
wire csrbank16_ev_pending_r;
reg csrbank16_ev_pending_we = 1'd0;
wire csrbank16_ev_pending_w;
reg csrbank16_ev_enable0_re = 1'd0;
wire csrbank16_ev_enable0_r;
reg csrbank16_ev_enable0_we = 1'd0;
wire csrbank16_ev_enable0_w;
wire csrbank16_sel;
wire [13:0] interface17_bank_bus_adr;
wire interface17_bank_bus_we;
wire [31:0] interface17_bank_bus_dat_w;
reg [31:0] interface17_bank_bus_dat_r = 32'd0;
reg csrbank17_in_re = 1'd0;
wire csrbank17_in_r;
reg csrbank17_in_we = 1'd0;
wire csrbank17_in_w;
reg csrbank17_mode0_re = 1'd0;
wire csrbank17_mode0_r;
reg csrbank17_mode0_we = 1'd0;
wire csrbank17_mode0_w;
reg csrbank17_edge0_re = 1'd0;
wire csrbank17_edge0_r;
reg csrbank17_edge0_we = 1'd0;
wire csrbank17_edge0_w;
reg csrbank17_ev_status_re = 1'd0;
wire csrbank17_ev_status_r;
reg csrbank17_ev_status_we = 1'd0;
wire csrbank17_ev_status_w;
reg csrbank17_ev_pending_re = 1'd0;
wire csrbank17_ev_pending_r;
reg csrbank17_ev_pending_we = 1'd0;
wire csrbank17_ev_pending_w;
reg csrbank17_ev_enable0_re = 1'd0;
wire csrbank17_ev_enable0_r;
reg csrbank17_ev_enable0_we = 1'd0;
wire csrbank17_ev_enable0_w;
wire csrbank17_sel;
wire [13:0] interface18_bank_bus_adr;
wire interface18_bank_bus_we;
wire [31:0] interface18_bank_bus_dat_w;
reg [31:0] interface18_bank_bus_dat_r = 32'd0;
reg csrbank18_in_re = 1'd0;
wire csrbank18_in_r;
reg csrbank18_in_we = 1'd0;
wire csrbank18_in_w;
reg csrbank18_mode0_re = 1'd0;
wire csrbank18_mode0_r;
reg csrbank18_mode0_we = 1'd0;
wire csrbank18_mode0_w;
reg csrbank18_edge0_re = 1'd0;
wire csrbank18_edge0_r;
reg csrbank18_edge0_we = 1'd0;
wire csrbank18_edge0_w;
reg csrbank18_ev_status_re = 1'd0;
wire csrbank18_ev_status_r;
reg csrbank18_ev_status_we = 1'd0;
wire csrbank18_ev_status_w;
reg csrbank18_ev_pending_re = 1'd0;
wire csrbank18_ev_pending_r;
reg csrbank18_ev_pending_we = 1'd0;
wire csrbank18_ev_pending_w;
reg csrbank18_ev_enable0_re = 1'd0;
wire csrbank18_ev_enable0_r;
reg csrbank18_ev_enable0_we = 1'd0;
wire csrbank18_ev_enable0_w;
wire csrbank18_sel;
wire [13:0] interface19_bank_bus_adr;
wire interface19_bank_bus_we;
wire [31:0] interface19_bank_bus_dat_w;
reg [31:0] interface19_bank_bus_dat_r = 32'd0;
reg csrbank19_out0_re = 1'd0;
wire [2:0] csrbank19_out0_r;
reg csrbank19_out0_we = 1'd0;
wire [2:0] csrbank19_out0_w;
wire csrbank19_sel;
wire [13:0] csr_interconnect_adr;
wire csr_interconnect_we;
wire [31:0] csr_interconnect_dat_w;
wire [31:0] csr_interconnect_dat_r;
reg state = 1'd0;
reg next_state = 1'd0;
reg [29:0] comb_array_muxed0 = 30'd0;
reg [31:0] comb_array_muxed1 = 32'd0;
reg [3:0] comb_array_muxed2 = 4'd0;
reg comb_array_muxed3 = 1'd0;
reg comb_array_muxed4 = 1'd0;
reg comb_array_muxed5 = 1'd0;
reg [2:0] comb_array_muxed6 = 3'd0;
reg [1:0] comb_array_muxed7 = 2'd0;
reg sync_array_muxed = 1'd0;
wire sdrio_clk;
wire sdrio_clk_1;
wire sdrio_clk_2;
wire sdrio_clk_3;
reg multiregimpl0_regs0 = 1'd0;
reg multiregimpl0_regs1 = 1'd0;
reg multiregimpl1_regs0 = 1'd0;
reg multiregimpl1_regs1 = 1'd0;
reg multiregimpl2_regs0 = 1'd0;
reg multiregimpl2_regs1 = 1'd0;
reg multiregimpl3_regs0 = 1'd0;
reg multiregimpl3_regs1 = 1'd0;
reg multiregimpl4_regs0 = 1'd0;
reg multiregimpl4_regs1 = 1'd0;
reg multiregimpl5_regs0 = 1'd0;
reg multiregimpl5_regs1 = 1'd0;
reg multiregimpl6_regs0 = 1'd0;
reg multiregimpl6_regs1 = 1'd0;
reg multiregimpl7_regs0 = 1'd0;
reg multiregimpl7_regs1 = 1'd0;
reg multiregimpl8_regs0 = 1'd0;
reg multiregimpl8_regs1 = 1'd0;
reg multiregimpl9_regs0 = 1'd0;
reg multiregimpl9_regs1 = 1'd0;
reg multiregimpl10_regs0 = 1'd0;
reg multiregimpl10_regs1 = 1'd0;
reg multiregimpl11_regs0 = 1'd0;
reg multiregimpl11_regs1 = 1'd0;
reg multiregimpl12_regs0 = 1'd0;
reg multiregimpl12_regs1 = 1'd0;
reg multiregimpl13_regs0 = 1'd0;
reg multiregimpl13_regs1 = 1'd0;
reg multiregimpl14_regs0 = 1'd0;
reg multiregimpl14_regs1 = 1'd0;
reg multiregimpl15_regs0 = 1'd0;
reg multiregimpl15_regs1 = 1'd0;
reg multiregimpl16_regs0 = 1'd0;
reg multiregimpl16_regs1 = 1'd0;
reg multiregimpl17_regs0 = 1'd0;
reg multiregimpl17_regs1 = 1'd0;
reg multiregimpl18_regs0 = 1'd0;
reg multiregimpl18_regs1 = 1'd0;
reg multiregimpl19_regs0 = 1'd0;
reg multiregimpl19_regs1 = 1'd0;
reg multiregimpl20_regs0 = 1'd0;
reg multiregimpl20_regs1 = 1'd0;
reg multiregimpl21_regs0 = 1'd0;
reg multiregimpl21_regs1 = 1'd0;
reg multiregimpl22_regs0 = 1'd0;
reg multiregimpl22_regs1 = 1'd0;
reg multiregimpl23_regs0 = 1'd0;
reg multiregimpl23_regs1 = 1'd0;
reg multiregimpl24_regs0 = 1'd0;
reg multiregimpl24_regs1 = 1'd0;
reg multiregimpl25_regs0 = 1'd0;
reg multiregimpl25_regs1 = 1'd0;
reg multiregimpl26_regs0 = 1'd0;
reg multiregimpl26_regs1 = 1'd0;
reg multiregimpl27_regs0 = 1'd0;
reg multiregimpl27_regs1 = 1'd0;
reg multiregimpl28_regs0 = 1'd0;
reg multiregimpl28_regs1 = 1'd0;
reg multiregimpl29_regs0 = 1'd0;
reg multiregimpl29_regs1 = 1'd0;
reg multiregimpl30_regs0 = 1'd0;
reg multiregimpl30_regs1 = 1'd0;
reg multiregimpl31_regs0 = 1'd0;
reg multiregimpl31_regs1 = 1'd0;
reg multiregimpl32_regs0 = 1'd0;
reg multiregimpl32_regs1 = 1'd0;
reg multiregimpl33_regs0 = 1'd0;
reg multiregimpl33_regs1 = 1'd0;
reg multiregimpl34_regs0 = 1'd0;
reg multiregimpl34_regs1 = 1'd0;
reg multiregimpl35_regs0 = 1'd0;
reg multiregimpl35_regs1 = 1'd0;
reg multiregimpl36_regs0 = 1'd0;
reg multiregimpl36_regs1 = 1'd0;
reg multiregimpl37_regs0 = 1'd0;
reg multiregimpl37_regs1 = 1'd0;
reg multiregimpl38_regs0 = 1'd0;
reg multiregimpl38_regs1 = 1'd0;
reg multiregimpl39_regs0 = 1'd0;
reg multiregimpl39_regs1 = 1'd0;
reg multiregimpl40_regs0 = 1'd0;
reg multiregimpl40_regs1 = 1'd0;
reg multiregimpl41_regs0 = 1'd0;
reg multiregimpl41_regs1 = 1'd0;
reg multiregimpl42_regs0 = 1'd0;
reg multiregimpl42_regs1 = 1'd0;
reg multiregimpl43_regs0 = 1'd0;
reg multiregimpl43_regs1 = 1'd0;
reg multiregimpl44_regs0 = 1'd0;
reg multiregimpl44_regs1 = 1'd0;
reg multiregimpl45_regs0 = 1'd0;
reg multiregimpl45_regs1 = 1'd0;
reg multiregimpl46_regs0 = 1'd0;
reg multiregimpl46_regs1 = 1'd0;
reg multiregimpl47_regs0 = 1'd0;
reg multiregimpl47_regs1 = 1'd0;
reg multiregimpl48_regs0 = 1'd0;
reg multiregimpl48_regs1 = 1'd0;
reg multiregimpl49_regs0 = 1'd0;
reg multiregimpl49_regs1 = 1'd0;
reg multiregimpl50_regs0 = 1'd0;
reg multiregimpl50_regs1 = 1'd0;
reg multiregimpl51_regs0 = 1'd0;
reg multiregimpl51_regs1 = 1'd0;
reg multiregimpl52_regs0 = 1'd0;
reg multiregimpl52_regs1 = 1'd0;
reg multiregimpl53_regs0 = 1'd0;
reg multiregimpl53_regs1 = 1'd0;
reg multiregimpl54_regs0 = 1'd0;
reg multiregimpl54_regs1 = 1'd0;
reg multiregimpl55_regs0 = 1'd0;
reg multiregimpl55_regs1 = 1'd0;
reg multiregimpl56_regs0 = 1'd0;
reg multiregimpl56_regs1 = 1'd0;
reg multiregimpl57_regs0 = 1'd0;
reg multiregimpl57_regs1 = 1'd0;
reg multiregimpl58_regs0 = 1'd0;
reg multiregimpl58_regs1 = 1'd0;
reg multiregimpl59_regs0 = 1'd0;
reg multiregimpl59_regs1 = 1'd0;
reg multiregimpl60_regs0 = 1'd0;
reg multiregimpl60_regs1 = 1'd0;
reg multiregimpl61_regs0 = 1'd0;
reg multiregimpl61_regs1 = 1'd0;
reg multiregimpl62_regs0 = 1'd0;
reg multiregimpl62_regs1 = 1'd0;
reg multiregimpl63_regs0 = 1'd0;
reg multiregimpl63_regs1 = 1'd0;
reg multiregimpl64_regs0 = 1'd0;
reg multiregimpl64_regs1 = 1'd0;
reg multiregimpl65_regs0 = 1'd0;
reg multiregimpl65_regs1 = 1'd0;
reg multiregimpl66_regs0 = 1'd0;
reg multiregimpl66_regs1 = 1'd0;
reg multiregimpl67_regs0 = 1'd0;
reg multiregimpl67_regs1 = 1'd0;
reg multiregimpl68_regs0 = 1'd0;
reg multiregimpl68_regs1 = 1'd0;
reg multiregimpl69_regs0 = 1'd0;
reg multiregimpl69_regs1 = 1'd0;
reg multiregimpl70_regs0 = 1'd0;
reg multiregimpl70_regs1 = 1'd0;
reg multiregimpl71_regs0 = 1'd0;
reg multiregimpl71_regs1 = 1'd0;
reg multiregimpl72_regs0 = 1'd0;
reg multiregimpl72_regs1 = 1'd0;
reg multiregimpl73_regs0 = 1'd0;
reg multiregimpl73_regs1 = 1'd0;
reg multiregimpl74_regs0 = 1'd0;
reg multiregimpl74_regs1 = 1'd0;
reg multiregimpl75_regs0 = 1'd0;
reg multiregimpl75_regs1 = 1'd0;
reg multiregimpl76_regs0 = 1'd0;
reg multiregimpl76_regs1 = 1'd0;
reg multiregimpl77_regs0 = 1'd0;
reg multiregimpl77_regs1 = 1'd0;
reg multiregimpl78_regs0 = 1'd0;
reg multiregimpl78_regs1 = 1'd0;
reg multiregimpl79_regs0 = 1'd0;
reg multiregimpl79_regs1 = 1'd0;
reg multiregimpl80_regs0 = 1'd0;
reg multiregimpl80_regs1 = 1'd0;
reg multiregimpl81_regs0 = 1'd0;
reg multiregimpl81_regs1 = 1'd0;
reg multiregimpl82_regs0 = 1'd0;
reg multiregimpl82_regs1 = 1'd0;
reg multiregimpl83_regs0 = 1'd0;
reg multiregimpl83_regs1 = 1'd0;
reg multiregimpl84_regs0 = 1'd0;
reg multiregimpl84_regs1 = 1'd0;
reg multiregimpl85_regs0 = 1'd0;
reg multiregimpl85_regs1 = 1'd0;
reg multiregimpl86_regs0 = 1'd0;
reg multiregimpl86_regs1 = 1'd0;
reg multiregimpl87_regs0 = 1'd0;
reg multiregimpl87_regs1 = 1'd0;
reg multiregimpl88_regs0 = 1'd0;
reg multiregimpl88_regs1 = 1'd0;
reg multiregimpl89_regs0 = 1'd0;
reg multiregimpl89_regs1 = 1'd0;
reg multiregimpl90_regs0 = 1'd0;
reg multiregimpl90_regs1 = 1'd0;
reg multiregimpl91_regs0 = 1'd0;
reg multiregimpl91_regs1 = 1'd0;
reg multiregimpl92_regs0 = 1'd0;
reg multiregimpl92_regs1 = 1'd0;
reg multiregimpl93_regs0 = 1'd0;
reg multiregimpl93_regs1 = 1'd0;
reg multiregimpl94_regs0 = 1'd0;
reg multiregimpl94_regs1 = 1'd0;
reg multiregimpl95_regs0 = 1'd0;
reg multiregimpl95_regs1 = 1'd0;
reg multiregimpl96_regs0 = 1'd0;
reg multiregimpl96_regs1 = 1'd0;
reg multiregimpl97_regs0 = 1'd0;
reg multiregimpl97_regs1 = 1'd0;
reg multiregimpl98_regs0 = 1'd0;
reg multiregimpl98_regs1 = 1'd0;
reg multiregimpl99_regs0 = 1'd0;
reg multiregimpl99_regs1 = 1'd0;
reg multiregimpl100_regs0 = 1'd0;
reg multiregimpl100_regs1 = 1'd0;
reg multiregimpl101_regs0 = 1'd0;
reg multiregimpl101_regs1 = 1'd0;
reg multiregimpl102_regs0 = 1'd0;
reg multiregimpl102_regs1 = 1'd0;
reg multiregimpl103_regs0 = 1'd0;
reg multiregimpl103_regs1 = 1'd0;
reg multiregimpl104_regs0 = 1'd0;
reg multiregimpl104_regs1 = 1'd0;
reg multiregimpl105_regs0 = 1'd0;
reg multiregimpl105_regs1 = 1'd0;
reg multiregimpl106_regs0 = 1'd0;
reg multiregimpl106_regs1 = 1'd0;
reg multiregimpl107_regs0 = 1'd0;
reg multiregimpl107_regs1 = 1'd0;
reg multiregimpl108_regs0 = 1'd0;
reg multiregimpl108_regs1 = 1'd0;
reg multiregimpl109_regs0 = 1'd0;
reg multiregimpl109_regs1 = 1'd0;
reg multiregimpl110_regs0 = 1'd0;
reg multiregimpl110_regs1 = 1'd0;
reg multiregimpl111_regs0 = 1'd0;
reg multiregimpl111_regs1 = 1'd0;
reg multiregimpl112_regs0 = 1'd0;
reg multiregimpl112_regs1 = 1'd0;
reg multiregimpl113_regs0 = 1'd0;
reg multiregimpl113_regs1 = 1'd0;
reg multiregimpl114_regs0 = 1'd0;
reg multiregimpl114_regs1 = 1'd0;
reg multiregimpl115_regs0 = 1'd0;
reg multiregimpl115_regs1 = 1'd0;
reg multiregimpl116_regs0 = 1'd0;
reg multiregimpl116_regs1 = 1'd0;
reg multiregimpl117_regs0 = 1'd0;
reg multiregimpl117_regs1 = 1'd0;
reg multiregimpl118_regs0 = 1'd0;
reg multiregimpl118_regs1 = 1'd0;
reg multiregimpl119_regs0 = 1'd0;
reg multiregimpl119_regs1 = 1'd0;
reg multiregimpl120_regs0 = 1'd0;
reg multiregimpl120_regs1 = 1'd0;
reg multiregimpl121_regs0 = 1'd0;
reg multiregimpl121_regs1 = 1'd0;
reg multiregimpl122_regs0 = 1'd0;
reg multiregimpl122_regs1 = 1'd0;
reg multiregimpl123_regs0 = 1'd0;
reg multiregimpl123_regs1 = 1'd0;
reg multiregimpl124_regs0 = 1'd0;
reg multiregimpl124_regs1 = 1'd0;
reg multiregimpl125_regs0 = 1'd0;
reg multiregimpl125_regs1 = 1'd0;
reg multiregimpl126_regs0 = 1'd0;
reg multiregimpl126_regs1 = 1'd0;
reg multiregimpl127_regs0 = 1'd0;
reg multiregimpl127_regs1 = 1'd0;
reg multiregimpl128_regs0 = 1'd0;
reg multiregimpl128_regs1 = 1'd0;
reg multiregimpl129_regs0 = 1'd0;
reg multiregimpl129_regs1 = 1'd0;
reg multiregimpl130_regs0 = 1'd0;
reg multiregimpl130_regs1 = 1'd0;
reg multiregimpl131_regs0 = 1'd0;
reg multiregimpl131_regs1 = 1'd0;
reg multiregimpl132_regs0 = 1'd0;
reg multiregimpl132_regs1 = 1'd0;
reg multiregimpl133_regs0 = 1'd0;
reg multiregimpl133_regs1 = 1'd0;
reg multiregimpl134_regs0 = 1'd0;
reg multiregimpl134_regs1 = 1'd0;
reg multiregimpl135_regs0 = 1'd0;
reg multiregimpl135_regs1 = 1'd0;
reg multiregimpl136_regs0 = 1'd0;
reg multiregimpl136_regs1 = 1'd0;

assign core_rst = (~core_rstn);
assign mgmtsoc_reset = (mgmtsoc_soc_rst | mgmtsoc_cpu_rst);
assign spi_sdoenb = (~spi_cs_n);
assign mprj_cyc_o = mprj_cyc;
assign mprj_stb_o = mprj_stb;
assign mprj_we_o = mprj_we;
assign mprj_sel_o = mprj_sel;
always @(*) begin
	mprj_adr_o = 32'd0;
	mprj_adr_o[31:2] = mprj_adr;
	mprj_adr_o[1:0] = 1'd0;
end
assign mprj_dat_r = mprj_dat_i;
assign mprj_dat_o = mprj_dat_w;
assign mprj_ack = mprj_ack_i;
assign hk_stb_o = hk_stb;
assign hk_cyc_o = hk_cyc;
assign hk_dat_r = hk_dat_i;
assign hk_ack = hk_ack_i;
assign debug_out = 1'd0;
always @(*) begin
	sys_uart_rx = 1'd0;
	if ((debug_in == 1'd1)) begin
	end else begin
		sys_uart_rx = serial_rx;
	end
end
always @(*) begin
	dbg_uart_dbg_uart_rx = 1'd0;
	if ((debug_in == 1'd1)) begin
		dbg_uart_dbg_uart_rx = serial_rx;
	end else begin
	end
end
always @(*) begin
	serial_tx = 1'd0;
	if ((debug_in == 1'd1)) begin
		serial_tx = dbg_uart_dbg_uart_tx;
	end else begin
		serial_tx = sys_uart_tx;
	end
end
assign uart_enabled = (uart_enabled_o | debug_in);
assign qspi_enabled = 1'd0;
assign trap = 1'd0;
assign clk_out = clk_in;
assign resetn_out = resetn_in;
assign serial_load_out = serial_load_in;
assign serial_data_2_out = serial_data_2_in;
assign serial_resetn_out = serial_resetn_in;
assign serial_clock_out = serial_clock_in;
assign rstb_l_out = rstb_l_in;
assign por_l_out = por_l_in;
assign porb_h_out = porb_h_in;
assign mgmtsoc_bus_error = error;
always @(*) begin
	mgmtsoc_interrupt = 32'd0;
	mgmtsoc_interrupt[0] = mgmtsoc_irq;
	mgmtsoc_interrupt[1] = uart_irq;
	mgmtsoc_interrupt[2] = gpioin0_gpioin0_irq;
	mgmtsoc_interrupt[3] = gpioin1_gpioin1_irq;
	mgmtsoc_interrupt[4] = gpioin2_gpioin2_irq;
	mgmtsoc_interrupt[5] = gpioin3_gpioin3_irq;
	mgmtsoc_interrupt[6] = gpioin4_gpioin4_irq;
	mgmtsoc_interrupt[7] = gpioin5_gpioin5_irq;
end
assign sys_clk = core_clk;
assign por_clk = core_clk;
assign sys_rst = int_rst;
assign mgmtsoc_bus_errors_status = mgmtsoc_bus_errors;
assign mgmtsoc_zero_trigger = (mgmtsoc_value == 1'd0);
assign mgmtsoc_zero0 = mgmtsoc_zero_status;
assign mgmtsoc_zero1 = mgmtsoc_zero_pending;
always @(*) begin
	mgmtsoc_zero_clear = 1'd0;
	if ((mgmtsoc_pending_re & mgmtsoc_pending_r)) begin
		mgmtsoc_zero_clear = 1'd1;
	end
end
assign mgmtsoc_irq = (mgmtsoc_pending_status & mgmtsoc_enable_storage);
assign mgmtsoc_zero_status = mgmtsoc_zero_trigger;
assign dff_di = dff_bus_dat_w[31:0];
always @(*) begin
	dff_we = 4'd0;
	dff_we[0] = (((dff_bus_sel[0] & dff_bus_we) & dff_bus_stb) & dff_bus_cyc);
	dff_we[1] = (((dff_bus_sel[1] & dff_bus_we) & dff_bus_stb) & dff_bus_cyc);
	dff_we[2] = (((dff_bus_sel[2] & dff_bus_we) & dff_bus_stb) & dff_bus_cyc);
	dff_we[3] = (((dff_bus_sel[3] & dff_bus_we) & dff_bus_stb) & dff_bus_cyc);
end
assign dff_bus_dat_r[31:0] = dff_do;
assign dff_en = (dff_bus_stb & dff_bus_cyc);
assign dff2_di = dff2_bus_dat_w[31:0];
always @(*) begin
	dff2_we = 4'd0;
	dff2_we[0] = (((dff2_bus_sel[0] & dff2_bus_we) & dff2_bus_stb) & dff2_bus_cyc);
	dff2_we[1] = (((dff2_bus_sel[1] & dff2_bus_we) & dff2_bus_stb) & dff2_bus_cyc);
	dff2_we[2] = (((dff2_bus_sel[2] & dff2_bus_we) & dff2_bus_stb) & dff2_bus_cyc);
	dff2_we[3] = (((dff2_bus_sel[3] & dff2_bus_we) & dff2_bus_stb) & dff2_bus_cyc);
end
assign dff2_bus_dat_r[31:0] = dff2_do;
assign dff2_en = (dff2_bus_stb & dff2_bus_cyc);
assign mgmtsoc_litespisdrphycore_div = mgmtsoc_litespisdrphycore_spi_clk_divisor;
assign mgmtsoc_litespisdrphycore_sample_cnt = 1'd1;
assign mgmtsoc_litespisdrphycore_update_cnt = 1'd1;
assign mgmtsoc_litespisdrphycore_wait = mgmtsoc_litespisdrphycore_cs;
assign mgmtsoc_litespisdrphycore_cs_enable = mgmtsoc_litespisdrphycore_done;
assign flash_cs_n = (~mgmtsoc_litespisdrphycore_cs_enable);
assign flash_io1_oeb = 1'd1;
assign flash_io1_do = 1'd0;
assign flash_io2_do = 1'd0;
assign flash_io3_do = 1'd0;
assign flash_io2_oeb = 1'd1;
assign flash_io3_oeb = 1'd1;
assign mgmtsoc_litespisdrphycore_dq_oe = mgmtsoc_litespisdrphycore_sink_payload_mask;
always @(*) begin
	mgmtsoc_litespisdrphycore_dq_o = 1'd0;
	case (mgmtsoc_litespisdrphycore_sink_payload_width)
		1'd1: begin
			mgmtsoc_litespisdrphycore_dq_o = mgmtsoc_litespisdrphycore_sr_out[31];
		end
		2'd2: begin
			mgmtsoc_litespisdrphycore_dq_o = mgmtsoc_litespisdrphycore_sr_out[31:30];
		end
		3'd4: begin
			mgmtsoc_litespisdrphycore_dq_o = mgmtsoc_litespisdrphycore_sr_out[31:28];
		end
		4'd8: begin
			mgmtsoc_litespisdrphycore_dq_o = mgmtsoc_litespisdrphycore_sr_out[31:24];
		end
	endcase
end
assign mgmtsoc_litespisdrphycore_source_payload_data = mgmtsoc_litespisdrphycore_sr_in;
assign mgmtsoc_litespisdrphycore_spi_clk_divisor = mgmtsoc_litespisdrphycore_storage;
assign mgmtsoc_litespisdrphycore_posedge = ((mgmtsoc_litespisdrphycore_en & (~mgmtsoc_litespisdrphycore_clk)) & (mgmtsoc_litespisdrphycore_cnt == mgmtsoc_litespisdrphycore_div));
assign mgmtsoc_litespisdrphycore_negedge = ((mgmtsoc_litespisdrphycore_en & mgmtsoc_litespisdrphycore_clk) & (mgmtsoc_litespisdrphycore_cnt == mgmtsoc_litespisdrphycore_div));
assign mgmtsoc_litespisdrphycore_sample = (mgmtsoc_litespisdrphycore_cnt == mgmtsoc_litespisdrphycore_sample_cnt);
assign mgmtsoc_litespisdrphycore_update = (mgmtsoc_litespisdrphycore_cnt == mgmtsoc_litespisdrphycore_update_cnt);
assign mgmtsoc_litespisdrphycore_done = (mgmtsoc_litespisdrphycore_count == 1'd0);
always @(*) begin
	litespiphy_next_state = 2'd0;
	litespiphy_next_state = litespiphy_state;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_negedge) begin
				if ((mgmtsoc_litespisdrphycore_sr_cnt == 1'd0)) begin
					litespiphy_next_state = 2'd2;
				end
			end
		end
		2'd2: begin
			if (((mgmtsoc_litespisdrphycore_spi_clk_divisor > 1'd0) | mgmtsoc_litespisdrphycore_posedge_reg2)) begin
				litespiphy_next_state = 2'd3;
			end
		end
		2'd3: begin
			if (mgmtsoc_litespisdrphycore_source_ready) begin
				litespiphy_next_state = 1'd0;
			end
		end
		default: begin
			if ((mgmtsoc_litespisdrphycore_cs_enable & mgmtsoc_litespisdrphycore_sink_valid)) begin
				litespiphy_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sink_ready = 1'd0;
	case (litespiphy_state)
		1'd1: begin
		end
		2'd2: begin
			if (((mgmtsoc_litespisdrphycore_spi_clk_divisor > 1'd0) | mgmtsoc_litespisdrphycore_posedge_reg2)) begin
				mgmtsoc_litespisdrphycore_sink_ready = 1'd1;
			end
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_en = 1'd0;
	case (litespiphy_state)
		1'd1: begin
			mgmtsoc_litespisdrphycore_en = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value = 8'd0;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_negedge) begin
				mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value = (mgmtsoc_litespisdrphycore_sr_cnt - mgmtsoc_litespisdrphycore_sink_payload_width);
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			if ((mgmtsoc_litespisdrphycore_cs_enable & mgmtsoc_litespisdrphycore_sink_valid)) begin
				mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value = (mgmtsoc_litespisdrphycore_sink_payload_len - mgmtsoc_litespisdrphycore_sink_payload_width);
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_out_load = 1'd0;
	case (litespiphy_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			if ((mgmtsoc_litespisdrphycore_cs_enable & mgmtsoc_litespisdrphycore_sink_valid)) begin
				mgmtsoc_litespisdrphycore_sr_out_load = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce = 1'd0;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_negedge) begin
				mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce = 1'd1;
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			if ((mgmtsoc_litespisdrphycore_cs_enable & mgmtsoc_litespisdrphycore_sink_valid)) begin
				mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_out_shift = 1'd0;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_negedge) begin
				mgmtsoc_litespisdrphycore_sr_out_shift = 1'd1;
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_sr_in_shift = 1'd0;
	case (litespiphy_state)
		1'd1: begin
			if (mgmtsoc_litespisdrphycore_posedge_reg2) begin
				mgmtsoc_litespisdrphycore_sr_in_shift = 1'd1;
			end
		end
		2'd2: begin
			if (((mgmtsoc_litespisdrphycore_spi_clk_divisor > 1'd0) | mgmtsoc_litespisdrphycore_posedge_reg2)) begin
				mgmtsoc_litespisdrphycore_sr_in_shift = (mgmtsoc_litespisdrphycore_spi_clk_divisor == 1'd0);
			end
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_source_valid = 1'd0;
	case (litespiphy_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespisdrphycore_source_valid = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespisdrphycore_source_last = 1'd0;
	case (litespiphy_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespisdrphycore_source_last = 1'd1;
		end
		default: begin
		end
	endcase
end
assign mgmtsoc_litespisdrphycore_cs = mgmtsoc_crossbar_cs;
assign mgmtsoc_litespimmap_sink_valid = mgmtsoc_port_mmap_user_port_source_valid;
assign mgmtsoc_port_mmap_user_port_source_ready = mgmtsoc_litespimmap_sink_ready;
assign mgmtsoc_litespimmap_sink_first = mgmtsoc_port_mmap_user_port_source_first;
assign mgmtsoc_litespimmap_sink_last = mgmtsoc_port_mmap_user_port_source_last;
assign mgmtsoc_litespimmap_sink_payload_data = mgmtsoc_port_mmap_user_port_source_payload_data;
assign mgmtsoc_port_mmap_user_port_sink_valid = mgmtsoc_litespimmap_source_valid;
assign mgmtsoc_litespimmap_source_ready = mgmtsoc_port_mmap_user_port_sink_ready;
assign mgmtsoc_port_mmap_user_port_sink_first = mgmtsoc_litespimmap_source_first;
assign mgmtsoc_port_mmap_user_port_sink_last = mgmtsoc_litespimmap_source_last;
assign mgmtsoc_port_mmap_user_port_sink_payload_data = mgmtsoc_litespimmap_source_payload_data;
assign mgmtsoc_port_mmap_user_port_sink_payload_len = mgmtsoc_litespimmap_source_payload_len;
assign mgmtsoc_port_mmap_user_port_sink_payload_width = mgmtsoc_litespimmap_source_payload_width;
assign mgmtsoc_port_mmap_user_port_sink_payload_mask = mgmtsoc_litespimmap_source_payload_mask;
assign mgmtsoc_master_sink_sink_valid = mgmtsoc_port_master_user_port_source_valid;
assign mgmtsoc_port_master_user_port_source_ready = mgmtsoc_master_sink_sink_ready;
assign mgmtsoc_master_sink_sink_first = mgmtsoc_port_master_user_port_source_first;
assign mgmtsoc_master_sink_sink_last = mgmtsoc_port_master_user_port_source_last;
assign mgmtsoc_master_sink_sink_payload_data = mgmtsoc_port_master_user_port_source_payload_data;
assign mgmtsoc_port_master_user_port_sink_valid = mgmtsoc_master_source_source_valid;
assign mgmtsoc_master_source_source_ready = mgmtsoc_port_master_user_port_sink_ready;
assign mgmtsoc_port_master_user_port_sink_first = mgmtsoc_master_source_source_first;
assign mgmtsoc_port_master_user_port_sink_last = mgmtsoc_master_source_source_last;
assign mgmtsoc_port_master_user_port_sink_payload_data = mgmtsoc_master_source_source_payload_data;
assign mgmtsoc_port_master_user_port_sink_payload_len = mgmtsoc_master_source_source_payload_len;
assign mgmtsoc_port_master_user_port_sink_payload_width = mgmtsoc_master_source_source_payload_width;
assign mgmtsoc_port_master_user_port_sink_payload_mask = mgmtsoc_master_source_source_payload_mask;
assign mgmtsoc_litespisdrphycore_sink_valid = mgmtsoc_crossbar_source_valid;
assign mgmtsoc_crossbar_source_ready = mgmtsoc_litespisdrphycore_sink_ready;
assign mgmtsoc_litespisdrphycore_sink_first = mgmtsoc_crossbar_source_first;
assign mgmtsoc_litespisdrphycore_sink_last = mgmtsoc_crossbar_source_last;
assign mgmtsoc_litespisdrphycore_sink_payload_data = mgmtsoc_crossbar_source_payload_data;
assign mgmtsoc_litespisdrphycore_sink_payload_len = mgmtsoc_crossbar_source_payload_len;
assign mgmtsoc_litespisdrphycore_sink_payload_width = mgmtsoc_crossbar_source_payload_width;
assign mgmtsoc_litespisdrphycore_sink_payload_mask = mgmtsoc_crossbar_source_payload_mask;
assign mgmtsoc_crossbar_sink_valid = mgmtsoc_litespisdrphycore_source_valid;
assign mgmtsoc_litespisdrphycore_source_ready = mgmtsoc_crossbar_sink_ready;
assign mgmtsoc_crossbar_sink_first = mgmtsoc_litespisdrphycore_source_first;
assign mgmtsoc_crossbar_sink_last = mgmtsoc_litespisdrphycore_source_last;
assign mgmtsoc_crossbar_sink_payload_data = mgmtsoc_litespisdrphycore_source_payload_data;
assign mgmtsoc_port_mmap_internal_port_sink_valid = mgmtsoc_port_mmap_user_port_sink_valid;
assign mgmtsoc_port_mmap_user_port_sink_ready = mgmtsoc_port_mmap_internal_port_sink_ready;
assign mgmtsoc_port_mmap_internal_port_sink_first = mgmtsoc_port_mmap_user_port_sink_first;
assign mgmtsoc_port_mmap_internal_port_sink_last = mgmtsoc_port_mmap_user_port_sink_last;
assign mgmtsoc_port_mmap_internal_port_sink_payload_data = mgmtsoc_port_mmap_user_port_sink_payload_data;
assign mgmtsoc_port_mmap_internal_port_sink_payload_len = mgmtsoc_port_mmap_user_port_sink_payload_len;
assign mgmtsoc_port_mmap_internal_port_sink_payload_width = mgmtsoc_port_mmap_user_port_sink_payload_width;
assign mgmtsoc_port_mmap_internal_port_sink_payload_mask = mgmtsoc_port_mmap_user_port_sink_payload_mask;
assign mgmtsoc_port_mmap_user_port_source_valid = mgmtsoc_port_mmap_internal_port_source_valid;
assign mgmtsoc_port_mmap_internal_port_source_ready = mgmtsoc_port_mmap_user_port_source_ready;
assign mgmtsoc_port_mmap_user_port_source_first = mgmtsoc_port_mmap_internal_port_source_first;
assign mgmtsoc_port_mmap_user_port_source_last = mgmtsoc_port_mmap_internal_port_source_last;
assign mgmtsoc_port_mmap_user_port_source_payload_data = mgmtsoc_port_mmap_internal_port_source_payload_data;
assign mgmtsoc_port_mmap_request = mgmtsoc_litespimmap_cs;
assign mgmtsoc_port_master_internal_port_sink_valid = mgmtsoc_port_master_user_port_sink_valid;
assign mgmtsoc_port_master_user_port_sink_ready = mgmtsoc_port_master_internal_port_sink_ready;
assign mgmtsoc_port_master_internal_port_sink_first = mgmtsoc_port_master_user_port_sink_first;
assign mgmtsoc_port_master_internal_port_sink_last = mgmtsoc_port_master_user_port_sink_last;
assign mgmtsoc_port_master_internal_port_sink_payload_data = mgmtsoc_port_master_user_port_sink_payload_data;
assign mgmtsoc_port_master_internal_port_sink_payload_len = mgmtsoc_port_master_user_port_sink_payload_len;
assign mgmtsoc_port_master_internal_port_sink_payload_width = mgmtsoc_port_master_user_port_sink_payload_width;
assign mgmtsoc_port_master_internal_port_sink_payload_mask = mgmtsoc_port_master_user_port_sink_payload_mask;
assign mgmtsoc_port_master_user_port_source_valid = mgmtsoc_port_master_internal_port_source_valid;
assign mgmtsoc_port_master_internal_port_source_ready = mgmtsoc_port_master_user_port_source_ready;
assign mgmtsoc_port_master_user_port_source_first = mgmtsoc_port_master_internal_port_source_first;
assign mgmtsoc_port_master_user_port_source_last = mgmtsoc_port_master_internal_port_source_last;
assign mgmtsoc_port_master_user_port_source_payload_data = mgmtsoc_port_master_internal_port_source_payload_data;
assign mgmtsoc_port_master_request = mgmtsoc_master_cs;
assign litespi_tx_mux_endpoint0_sink_valid = mgmtsoc_port_mmap_internal_port_sink_valid;
assign mgmtsoc_port_mmap_internal_port_sink_ready = litespi_tx_mux_endpoint0_sink_ready;
assign litespi_tx_mux_endpoint0_sink_first = mgmtsoc_port_mmap_internal_port_sink_first;
assign litespi_tx_mux_endpoint0_sink_last = mgmtsoc_port_mmap_internal_port_sink_last;
assign litespi_tx_mux_endpoint0_sink_payload_data = mgmtsoc_port_mmap_internal_port_sink_payload_data;
assign litespi_tx_mux_endpoint0_sink_payload_len = mgmtsoc_port_mmap_internal_port_sink_payload_len;
assign litespi_tx_mux_endpoint0_sink_payload_width = mgmtsoc_port_mmap_internal_port_sink_payload_width;
assign litespi_tx_mux_endpoint0_sink_payload_mask = mgmtsoc_port_mmap_internal_port_sink_payload_mask;
assign mgmtsoc_port_mmap_internal_port_source_valid = litespi_rx_demux_endpoint0_source_valid;
assign litespi_rx_demux_endpoint0_source_ready = mgmtsoc_port_mmap_internal_port_source_ready;
assign mgmtsoc_port_mmap_internal_port_source_first = litespi_rx_demux_endpoint0_source_first;
assign mgmtsoc_port_mmap_internal_port_source_last = litespi_rx_demux_endpoint0_source_last;
assign mgmtsoc_port_mmap_internal_port_source_payload_data = litespi_rx_demux_endpoint0_source_payload_data;
assign litespi_tx_mux_endpoint1_sink_valid = mgmtsoc_port_master_internal_port_sink_valid;
assign mgmtsoc_port_master_internal_port_sink_ready = litespi_tx_mux_endpoint1_sink_ready;
assign litespi_tx_mux_endpoint1_sink_first = mgmtsoc_port_master_internal_port_sink_first;
assign litespi_tx_mux_endpoint1_sink_last = mgmtsoc_port_master_internal_port_sink_last;
assign litespi_tx_mux_endpoint1_sink_payload_data = mgmtsoc_port_master_internal_port_sink_payload_data;
assign litespi_tx_mux_endpoint1_sink_payload_len = mgmtsoc_port_master_internal_port_sink_payload_len;
assign litespi_tx_mux_endpoint1_sink_payload_width = mgmtsoc_port_master_internal_port_sink_payload_width;
assign litespi_tx_mux_endpoint1_sink_payload_mask = mgmtsoc_port_master_internal_port_sink_payload_mask;
assign mgmtsoc_port_master_internal_port_source_valid = litespi_rx_demux_endpoint1_source_valid;
assign litespi_rx_demux_endpoint1_source_ready = mgmtsoc_port_master_internal_port_source_ready;
assign mgmtsoc_port_master_internal_port_source_first = litespi_rx_demux_endpoint1_source_first;
assign mgmtsoc_port_master_internal_port_source_last = litespi_rx_demux_endpoint1_source_last;
assign mgmtsoc_port_master_internal_port_source_payload_data = litespi_rx_demux_endpoint1_source_payload_data;
assign litespi_request = {mgmtsoc_port_master_request, mgmtsoc_port_mmap_request};
assign mgmtsoc_crossbar_source_valid = litespi_tx_mux_source_valid;
assign litespi_tx_mux_source_ready = mgmtsoc_crossbar_source_ready;
assign mgmtsoc_crossbar_source_first = litespi_tx_mux_source_first;
assign mgmtsoc_crossbar_source_last = litespi_tx_mux_source_last;
assign mgmtsoc_crossbar_source_payload_data = litespi_tx_mux_source_payload_data;
assign mgmtsoc_crossbar_source_payload_len = litespi_tx_mux_source_payload_len;
assign mgmtsoc_crossbar_source_payload_width = litespi_tx_mux_source_payload_width;
assign mgmtsoc_crossbar_source_payload_mask = litespi_tx_mux_source_payload_mask;
assign litespi_tx_mux_sel = litespi_grant;
assign litespi_rx_demux_sink_valid = mgmtsoc_crossbar_sink_valid;
assign mgmtsoc_crossbar_sink_ready = litespi_rx_demux_sink_ready;
assign litespi_rx_demux_sink_first = mgmtsoc_crossbar_sink_first;
assign litespi_rx_demux_sink_last = mgmtsoc_crossbar_sink_last;
assign litespi_rx_demux_sink_payload_data = mgmtsoc_crossbar_sink_payload_data;
assign litespi_rx_demux_sel = litespi_grant;
always @(*) begin
	mgmtsoc_crossbar_cs = 1'd0;
	case (litespi_grant)
		1'd0: begin
			mgmtsoc_crossbar_cs = mgmtsoc_litespimmap_cs;
		end
		1'd1: begin
			mgmtsoc_crossbar_cs = mgmtsoc_master_cs;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_valid = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_valid = litespi_tx_mux_endpoint0_sink_valid;
		end
		1'd1: begin
			litespi_tx_mux_source_valid = litespi_tx_mux_endpoint1_sink_valid;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_endpoint1_sink_ready = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_tx_mux_endpoint1_sink_ready = litespi_tx_mux_source_ready;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_first = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_first = litespi_tx_mux_endpoint0_sink_first;
		end
		1'd1: begin
			litespi_tx_mux_source_first = litespi_tx_mux_endpoint1_sink_first;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_last = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_last = litespi_tx_mux_endpoint0_sink_last;
		end
		1'd1: begin
			litespi_tx_mux_source_last = litespi_tx_mux_endpoint1_sink_last;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_payload_data = 32'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_payload_data = litespi_tx_mux_endpoint0_sink_payload_data;
		end
		1'd1: begin
			litespi_tx_mux_source_payload_data = litespi_tx_mux_endpoint1_sink_payload_data;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_payload_len = 6'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_payload_len = litespi_tx_mux_endpoint0_sink_payload_len;
		end
		1'd1: begin
			litespi_tx_mux_source_payload_len = litespi_tx_mux_endpoint1_sink_payload_len;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_payload_width = 4'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_payload_width = litespi_tx_mux_endpoint0_sink_payload_width;
		end
		1'd1: begin
			litespi_tx_mux_source_payload_width = litespi_tx_mux_endpoint1_sink_payload_width;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_source_payload_mask = 8'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_source_payload_mask = litespi_tx_mux_endpoint0_sink_payload_mask;
		end
		1'd1: begin
			litespi_tx_mux_source_payload_mask = litespi_tx_mux_endpoint1_sink_payload_mask;
		end
	endcase
end
always @(*) begin
	litespi_tx_mux_endpoint0_sink_ready = 1'd0;
	case (litespi_tx_mux_sel)
		1'd0: begin
			litespi_tx_mux_endpoint0_sink_ready = litespi_tx_mux_source_ready;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_sink_ready = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_sink_ready = litespi_rx_demux_endpoint0_source_ready;
		end
		1'd1: begin
			litespi_rx_demux_sink_ready = litespi_rx_demux_endpoint1_source_ready;
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint0_source_valid = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_endpoint0_source_valid = litespi_rx_demux_sink_valid;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint0_source_first = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_endpoint0_source_first = litespi_rx_demux_sink_first;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint0_source_last = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_endpoint0_source_last = litespi_rx_demux_sink_last;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint0_source_payload_data = 32'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
			litespi_rx_demux_endpoint0_source_payload_data = litespi_rx_demux_sink_payload_data;
		end
		1'd1: begin
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint1_source_valid = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_rx_demux_endpoint1_source_valid = litespi_rx_demux_sink_valid;
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint1_source_first = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_rx_demux_endpoint1_source_first = litespi_rx_demux_sink_first;
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint1_source_last = 1'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_rx_demux_endpoint1_source_last = litespi_rx_demux_sink_last;
		end
	endcase
end
always @(*) begin
	litespi_rx_demux_endpoint1_source_payload_data = 32'd0;
	case (litespi_rx_demux_sel)
		1'd0: begin
		end
		1'd1: begin
			litespi_rx_demux_endpoint1_source_payload_data = litespi_rx_demux_sink_payload_data;
		end
	endcase
end
assign mgmtsoc_litespimmap_spi_dummy_bits = mgmtsoc_litespimmap_storage;
assign mgmtsoc_litespimmap_done = (mgmtsoc_litespimmap_count == 1'd0);
always @(*) begin
	litespi_next_state = 4'd0;
	litespi_next_state = litespi_state;
	case (litespi_state)
		1'd1: begin
			if (mgmtsoc_litespimmap_source_ready) begin
				litespi_next_state = 2'd2;
			end
		end
		2'd2: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				litespi_next_state = 2'd3;
			end
		end
		2'd3: begin
			if (mgmtsoc_litespimmap_source_ready) begin
				litespi_next_state = 3'd4;
			end
		end
		3'd4: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				if ((mgmtsoc_litespimmap_spi_dummy_bits == 1'd0)) begin
					litespi_next_state = 3'd7;
				end else begin
					litespi_next_state = 3'd5;
				end
			end
		end
		3'd5: begin
			if (mgmtsoc_litespimmap_source_ready) begin
				litespi_next_state = 3'd6;
			end
		end
		3'd6: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				litespi_next_state = 3'd7;
			end
		end
		3'd7: begin
			if (mgmtsoc_litespimmap_source_ready) begin
				litespi_next_state = 4'd8;
			end
		end
		4'd8: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				litespi_next_state = 1'd0;
			end
		end
		default: begin
			if (((mgmtsoc_litespimmap_bus_cyc & mgmtsoc_litespimmap_bus_stb) & (~mgmtsoc_litespimmap_bus_we))) begin
				if ((mgmtsoc_litespimmap_burst_cs & (mgmtsoc_litespimmap_bus_adr == mgmtsoc_litespimmap_burst_adr))) begin
					litespi_next_state = 3'd7;
				end else begin
					litespi_next_state = 1'd1;
				end
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_bus_dat_r = 32'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
			mgmtsoc_litespimmap_bus_dat_r = {mgmtsoc_litespimmap_sink_payload_data[7:0], mgmtsoc_litespimmap_sink_payload_data[15:8], mgmtsoc_litespimmap_sink_payload_data[23:16], mgmtsoc_litespimmap_sink_payload_data[31:24]};
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_valid = 1'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_valid = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_valid = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_valid = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_valid = 1'd1;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
		end
		default: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value0 = (mgmtsoc_litespimmap_burst_cs & (~mgmtsoc_litespimmap_done));
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
		end
		default: begin
			mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_last = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_last = 1'd1;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_bus_ack = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				mgmtsoc_litespimmap_bus_ack = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_payload_data = 32'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_payload_data = 2'd3;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_payload_data = {mgmtsoc_litespimmap_bus_adr, mgmtsoc_litespimmap};
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_payload_data = mgmtsoc_litespimmap_dummy;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_payload_len = 6'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_payload_len = 4'd8;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_payload_len = 5'd24;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_payload_len = mgmtsoc_litespimmap_spi_dummy_bits;
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_payload_len = 6'd32;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_payload_width = 4'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_payload_width = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_payload_width = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_payload_width = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_payload_width = 1'd1;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_source_payload_mask = 8'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_source_payload_mask = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_source_payload_mask = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_source_payload_mask = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
			mgmtsoc_litespimmap_source_payload_mask = 1'd0;
		end
		4'd8: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = 30'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = mgmtsoc_litespimmap_bus_adr;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = mgmtsoc_litespimmap_bus_adr;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = mgmtsoc_litespimmap_bus_adr;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				mgmtsoc_litespimmap_burst_adr_litespi_next_value1 = (mgmtsoc_litespimmap_burst_adr + 1'd1);
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_cs = 1'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		2'd2: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		2'd3: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		3'd4: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		3'd5: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		3'd6: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		3'd7: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		4'd8: begin
			mgmtsoc_litespimmap_cs = 1'd1;
		end
		default: begin
			mgmtsoc_litespimmap_cs = mgmtsoc_litespimmap_burst_cs;
			if (((mgmtsoc_litespimmap_bus_cyc & mgmtsoc_litespimmap_bus_stb) & (~mgmtsoc_litespimmap_bus_we))) begin
				if ((mgmtsoc_litespimmap_burst_cs & (mgmtsoc_litespimmap_bus_adr == mgmtsoc_litespimmap_burst_adr))) begin
				end else begin
					mgmtsoc_litespimmap_cs = 1'd0;
				end
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd0;
	case (litespi_state)
		1'd1: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd1;
		end
		2'd2: begin
		end
		2'd3: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd1;
		end
		3'd4: begin
		end
		3'd5: begin
			mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd1;
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
			if (mgmtsoc_litespimmap_sink_valid) begin
				mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1 = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_sink_ready = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
			mgmtsoc_litespimmap_sink_ready = 1'd1;
		end
		2'd3: begin
		end
		3'd4: begin
			mgmtsoc_litespimmap_sink_ready = 1'd1;
		end
		3'd5: begin
		end
		3'd6: begin
			mgmtsoc_litespimmap_sink_ready = 1'd1;
		end
		3'd7: begin
		end
		4'd8: begin
			mgmtsoc_litespimmap_sink_ready = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_litespimmap_wait = 1'd0;
	case (litespi_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		3'd7: begin
		end
		4'd8: begin
		end
		default: begin
			mgmtsoc_litespimmap_wait = 1'd1;
		end
	endcase
end
assign mgmtsoc_master_rx_fifo_sink_valid = mgmtsoc_master_sink_sink_valid;
assign mgmtsoc_master_sink_sink_ready = mgmtsoc_master_rx_fifo_sink_ready;
assign mgmtsoc_master_rx_fifo_sink_first = mgmtsoc_master_sink_sink_first;
assign mgmtsoc_master_rx_fifo_sink_last = mgmtsoc_master_sink_sink_last;
assign mgmtsoc_master_rx_fifo_sink_payload_data = mgmtsoc_master_sink_sink_payload_data;
assign mgmtsoc_master_source_source_valid = mgmtsoc_master_tx_fifo_source_valid;
assign mgmtsoc_master_tx_fifo_source_ready = mgmtsoc_master_source_source_ready;
assign mgmtsoc_master_source_source_first = mgmtsoc_master_tx_fifo_source_first;
assign mgmtsoc_master_source_source_last = mgmtsoc_master_tx_fifo_source_last;
assign mgmtsoc_master_source_source_payload_data = mgmtsoc_master_tx_fifo_source_payload_data;
assign mgmtsoc_master_source_source_payload_len = mgmtsoc_master_tx_fifo_source_payload_len;
assign mgmtsoc_master_source_source_payload_width = mgmtsoc_master_tx_fifo_source_payload_width;
assign mgmtsoc_master_source_source_payload_mask = mgmtsoc_master_tx_fifo_source_payload_mask;
assign mgmtsoc_master_cs = mgmtsoc_master_cs_storage;
assign mgmtsoc_master_tx_fifo_sink_valid = mgmtsoc_master_rxtx_re;
assign mgmtsoc_master_tx_ready = mgmtsoc_master_tx_fifo_sink_ready;
assign mgmtsoc_master_tx_fifo_sink_payload_data = mgmtsoc_master_rxtx_r;
assign mgmtsoc_master_tx_fifo_sink_payload_len = mgmtsoc_master_len;
assign mgmtsoc_master_tx_fifo_sink_payload_width = mgmtsoc_master_width;
assign mgmtsoc_master_tx_fifo_sink_payload_mask = mgmtsoc_master_mask;
assign mgmtsoc_master_tx_fifo_sink_last = 1'd1;
assign mgmtsoc_master_rx_fifo_source_ready = mgmtsoc_master_rxtx_we;
assign mgmtsoc_master_rx_ready = mgmtsoc_master_rx_fifo_source_valid;
assign mgmtsoc_master_rxtx_w = mgmtsoc_master_rx_fifo_source_payload_data;
assign mgmtsoc_master_tx_fifo_sink_ready = ((~mgmtsoc_master_tx_fifo_source_valid) | mgmtsoc_master_tx_fifo_source_ready);
assign mgmtsoc_master_rx_fifo_sink_ready = ((~mgmtsoc_master_rx_fifo_source_valid) | mgmtsoc_master_rx_fifo_source_ready);
assign spi_master_start0 = spi_master_start1;
assign spi_master_length0 = spi_master_length1;
assign spi_master_done1 = spi_master_done0;
assign spi_master_mosi = spi_master_mosi_storage;
assign spi_master_miso_status = spi_master_miso;
assign spi_master_cs = spi_master_sel;
assign spi_master_cs_mode = spi_master_mode0;
assign spi_master_loopback = spi_master_mode1;
assign spi_master_clk_rise = (spi_master_clk_divider1 == (spi_master_clk_divider0[15:1] - 1'd1));
assign spi_master_clk_fall = (spi_master_clk_divider1 == (spi_master_clk_divider0 - 1'd1));
assign spi_master_clk_divider0 = spimaster_storage;
always @(*) begin
	spimaster_next_state = 2'd0;
	spimaster_next_state = spimaster_state;
	case (spimaster_state)
		1'd1: begin
			if (spi_master_clk_fall) begin
				spimaster_next_state = 2'd2;
			end
		end
		2'd2: begin
			if (spi_master_clk_fall) begin
				if ((spi_master_count == (spi_master_length0 - 1'd1))) begin
					spimaster_next_state = 2'd3;
				end
			end
		end
		2'd3: begin
			if (spi_master_clk_rise) begin
				spimaster_next_state = 1'd0;
			end
		end
		default: begin
			if (spi_master_start0) begin
				spimaster_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	spi_master_count_spimaster_next_value = 3'd0;
	case (spimaster_state)
		1'd1: begin
			spi_master_count_spimaster_next_value = 1'd0;
		end
		2'd2: begin
			if (spi_master_clk_fall) begin
				spi_master_count_spimaster_next_value = (spi_master_count + 1'd1);
			end
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_done0 = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			spi_master_done0 = 1'd1;
			if (spi_master_start0) begin
				spi_master_done0 = 1'd0;
			end
		end
	endcase
end
always @(*) begin
	spi_master_count_spimaster_next_value_ce = 1'd0;
	case (spimaster_state)
		1'd1: begin
			spi_master_count_spimaster_next_value_ce = 1'd1;
		end
		2'd2: begin
			if (spi_master_clk_fall) begin
				spi_master_count_spimaster_next_value_ce = 1'd1;
			end
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_irq = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			if (spi_master_clk_rise) begin
				spi_master_irq = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_clk_enable = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
			spi_master_clk_enable = 1'd1;
		end
		2'd3: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_xfer_enable = 1'd0;
	case (spimaster_state)
		1'd1: begin
			if (spi_master_clk_fall) begin
				spi_master_xfer_enable = 1'd1;
			end
		end
		2'd2: begin
			spi_master_xfer_enable = 1'd1;
		end
		2'd3: begin
			spi_master_xfer_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	spi_master_mosi_latch = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		default: begin
			if (spi_master_start0) begin
				spi_master_mosi_latch = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	spi_master_miso_latch = 1'd0;
	case (spimaster_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			if (spi_master_clk_rise) begin
				spi_master_miso_latch = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
assign mprj_wb_iena = mprj_wb_iena_storage;
always @(*) begin
	rs232phy_rs232phytx_next_state = 1'd0;
	rs232phy_rs232phytx_next_state = rs232phy_rs232phytx_state;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				if ((uart_phy_tx_count == 4'd9)) begin
					rs232phy_rs232phytx_next_state = 1'd0;
				end
			end
		end
		default: begin
			if (uart_phy_tx_sink_valid) begin
				rs232phy_rs232phytx_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd1;
			end
		end
		default: begin
			sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd1;
			if (uart_phy_tx_sink_valid) begin
				sys_uart_tx_rs232phy_rs232phytx_next_value_ce1 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	uart_phy_tx_data_rs232phy_rs232phytx_next_value2 = 8'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				uart_phy_tx_data_rs232phy_rs232phytx_next_value2 = {1'd1, uart_phy_tx_data[7:1]};
			end
		end
		default: begin
			if (uart_phy_tx_sink_valid) begin
				uart_phy_tx_data_rs232phy_rs232phytx_next_value2 = uart_phy_tx_sink_payload_data;
			end
		end
	endcase
end
always @(*) begin
	uart_phy_tx_sink_ready = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				if ((uart_phy_tx_count == 4'd9)) begin
					uart_phy_tx_sink_ready = 1'd1;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2 = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2 = 1'd1;
			end
		end
		default: begin
			if (uart_phy_tx_sink_valid) begin
				uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	uart_phy_tx_enable = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			uart_phy_tx_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_tx_count_rs232phy_rs232phytx_next_value0 = 4'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				uart_phy_tx_count_rs232phy_rs232phytx_next_value0 = (uart_phy_tx_count + 1'd1);
			end
		end
		default: begin
			uart_phy_tx_count_rs232phy_rs232phytx_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0 = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	sys_uart_tx_rs232phy_rs232phytx_next_value1 = 1'd0;
	case (rs232phy_rs232phytx_state)
		1'd1: begin
			if (uart_phy_tx_tick) begin
				sys_uart_tx_rs232phy_rs232phytx_next_value1 = uart_phy_tx_data;
			end
		end
		default: begin
			sys_uart_tx_rs232phy_rs232phytx_next_value1 = 1'd1;
			if (uart_phy_tx_sink_valid) begin
				sys_uart_tx_rs232phy_rs232phytx_next_value1 = 1'd0;
			end
		end
	endcase
end
always @(*) begin
	rs232phy_rs232phyrx_next_state = 1'd0;
	rs232phy_rs232phyrx_next_state = rs232phy_rs232phyrx_state;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				if ((uart_phy_rx_count == 4'd9)) begin
					rs232phy_rs232phyrx_next_state = 1'd0;
				end
			end
		end
		default: begin
			if (((uart_phy_rx_rx == 1'd0) & (uart_phy_rx_rx_d == 1'd1))) begin
				rs232phy_rs232phyrx_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	uart_phy_rx_data_rs232phy_rs232phyrx_next_value1 = 8'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				uart_phy_rx_data_rs232phy_rs232phyrx_next_value1 = {uart_phy_rx_rx, uart_phy_rx_data[7:1]};
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_data_rs232phy_rs232phyrx_next_value_ce1 = 1'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				uart_phy_rx_data_rs232phy_rs232phyrx_next_value_ce1 = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_source_valid = 1'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				if ((uart_phy_rx_count == 4'd9)) begin
					uart_phy_rx_source_valid = (uart_phy_rx_rx == 1'd1);
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_source_payload_data = 8'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				if ((uart_phy_rx_count == 4'd9)) begin
					uart_phy_rx_source_payload_data = uart_phy_rx_data;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_enable = 1'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			uart_phy_rx_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	uart_phy_rx_count_rs232phy_rs232phyrx_next_value0 = 4'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				uart_phy_rx_count_rs232phy_rs232phyrx_next_value0 = (uart_phy_rx_count + 1'd1);
			end
		end
		default: begin
			uart_phy_rx_count_rs232phy_rs232phyrx_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0 = 1'd0;
	case (rs232phy_rs232phyrx_state)
		1'd1: begin
			if (uart_phy_rx_tick) begin
				uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0 = 1'd1;
		end
	endcase
end
assign uart_uart_sink_valid = uart_phy_rx_source_valid;
assign uart_phy_rx_source_ready = uart_uart_sink_ready;
assign uart_uart_sink_first = uart_phy_rx_source_first;
assign uart_uart_sink_last = uart_phy_rx_source_last;
assign uart_uart_sink_payload_data = uart_phy_rx_source_payload_data;
assign uart_phy_tx_sink_valid = uart_uart_source_valid;
assign uart_uart_source_ready = uart_phy_tx_sink_ready;
assign uart_phy_tx_sink_first = uart_uart_source_first;
assign uart_phy_tx_sink_last = uart_uart_source_last;
assign uart_phy_tx_sink_payload_data = uart_uart_source_payload_data;
assign uart_tx_fifo_sink_valid = uart_rxtx_re;
assign uart_tx_fifo_sink_payload_data = uart_rxtx_r;
assign uart_uart_source_valid = uart_tx_fifo_source_valid;
assign uart_tx_fifo_source_ready = uart_uart_source_ready;
assign uart_uart_source_first = uart_tx_fifo_source_first;
assign uart_uart_source_last = uart_tx_fifo_source_last;
assign uart_uart_source_payload_data = uart_tx_fifo_source_payload_data;
assign uart_txfull_status = (~uart_tx_fifo_sink_ready);
assign uart_txempty_status = (~uart_tx_fifo_source_valid);
assign uart_tx_trigger = uart_tx_fifo_sink_ready;
assign uart_rx_fifo_sink_valid = uart_uart_sink_valid;
assign uart_uart_sink_ready = uart_rx_fifo_sink_ready;
assign uart_rx_fifo_sink_first = uart_uart_sink_first;
assign uart_rx_fifo_sink_last = uart_uart_sink_last;
assign uart_rx_fifo_sink_payload_data = uart_uart_sink_payload_data;
assign uart_rxtx_w = uart_rx_fifo_source_payload_data;
assign uart_rx_fifo_source_ready = (uart_rx_clear | (1'd0 & uart_rxtx_we));
assign uart_rxempty_status = (~uart_rx_fifo_source_valid);
assign uart_rxfull_status = (~uart_rx_fifo_sink_ready);
assign uart_rx_trigger = uart_rx_fifo_source_valid;
assign uart_tx0 = uart_tx_status;
assign uart_tx1 = uart_tx_pending;
always @(*) begin
	uart_tx_clear = 1'd0;
	if ((uart_pending_re & uart_pending_r[0])) begin
		uart_tx_clear = 1'd1;
	end
end
assign uart_rx0 = uart_rx_status;
assign uart_rx1 = uart_rx_pending;
always @(*) begin
	uart_rx_clear = 1'd0;
	if ((uart_pending_re & uart_pending_r[1])) begin
		uart_rx_clear = 1'd1;
	end
end
assign uart_irq = ((uart_pending_status[0] & uart_enable_storage[0]) | (uart_pending_status[1] & uart_enable_storage[1]));
assign uart_tx_status = uart_tx_trigger;
assign uart_rx_status = uart_rx_trigger;
assign uart_tx_fifo_syncfifo_din = {uart_tx_fifo_fifo_in_last, uart_tx_fifo_fifo_in_first, uart_tx_fifo_fifo_in_payload_data};
assign {uart_tx_fifo_fifo_out_last, uart_tx_fifo_fifo_out_first, uart_tx_fifo_fifo_out_payload_data} = uart_tx_fifo_syncfifo_dout;
assign uart_tx_fifo_sink_ready = uart_tx_fifo_syncfifo_writable;
assign uart_tx_fifo_syncfifo_we = uart_tx_fifo_sink_valid;
assign uart_tx_fifo_fifo_in_first = uart_tx_fifo_sink_first;
assign uart_tx_fifo_fifo_in_last = uart_tx_fifo_sink_last;
assign uart_tx_fifo_fifo_in_payload_data = uart_tx_fifo_sink_payload_data;
assign uart_tx_fifo_source_valid = uart_tx_fifo_readable;
assign uart_tx_fifo_source_first = uart_tx_fifo_fifo_out_first;
assign uart_tx_fifo_source_last = uart_tx_fifo_fifo_out_last;
assign uart_tx_fifo_source_payload_data = uart_tx_fifo_fifo_out_payload_data;
assign uart_tx_fifo_re = uart_tx_fifo_source_ready;
assign uart_tx_fifo_syncfifo_re = (uart_tx_fifo_syncfifo_readable & ((~uart_tx_fifo_readable) | uart_tx_fifo_re));
assign uart_tx_fifo_level1 = (uart_tx_fifo_level0 + uart_tx_fifo_readable);
always @(*) begin
	uart_tx_fifo_wrport_adr = 4'd0;
	if (uart_tx_fifo_replace) begin
		uart_tx_fifo_wrport_adr = (uart_tx_fifo_produce - 1'd1);
	end else begin
		uart_tx_fifo_wrport_adr = uart_tx_fifo_produce;
	end
end
assign uart_tx_fifo_wrport_dat_w = uart_tx_fifo_syncfifo_din;
assign uart_tx_fifo_wrport_we = (uart_tx_fifo_syncfifo_we & (uart_tx_fifo_syncfifo_writable | uart_tx_fifo_replace));
assign uart_tx_fifo_do_read = (uart_tx_fifo_syncfifo_readable & uart_tx_fifo_syncfifo_re);
assign uart_tx_fifo_rdport_adr = uart_tx_fifo_consume;
assign uart_tx_fifo_syncfifo_dout = uart_tx_fifo_rdport_dat_r;
assign uart_tx_fifo_rdport_re = uart_tx_fifo_do_read;
assign uart_tx_fifo_syncfifo_writable = (uart_tx_fifo_level0 != 5'd16);
assign uart_tx_fifo_syncfifo_readable = (uart_tx_fifo_level0 != 1'd0);
assign uart_rx_fifo_syncfifo_din = {uart_rx_fifo_fifo_in_last, uart_rx_fifo_fifo_in_first, uart_rx_fifo_fifo_in_payload_data};
assign {uart_rx_fifo_fifo_out_last, uart_rx_fifo_fifo_out_first, uart_rx_fifo_fifo_out_payload_data} = uart_rx_fifo_syncfifo_dout;
assign uart_rx_fifo_sink_ready = uart_rx_fifo_syncfifo_writable;
assign uart_rx_fifo_syncfifo_we = uart_rx_fifo_sink_valid;
assign uart_rx_fifo_fifo_in_first = uart_rx_fifo_sink_first;
assign uart_rx_fifo_fifo_in_last = uart_rx_fifo_sink_last;
assign uart_rx_fifo_fifo_in_payload_data = uart_rx_fifo_sink_payload_data;
assign uart_rx_fifo_source_valid = uart_rx_fifo_readable;
assign uart_rx_fifo_source_first = uart_rx_fifo_fifo_out_first;
assign uart_rx_fifo_source_last = uart_rx_fifo_fifo_out_last;
assign uart_rx_fifo_source_payload_data = uart_rx_fifo_fifo_out_payload_data;
assign uart_rx_fifo_re = uart_rx_fifo_source_ready;
assign uart_rx_fifo_syncfifo_re = (uart_rx_fifo_syncfifo_readable & ((~uart_rx_fifo_readable) | uart_rx_fifo_re));
assign uart_rx_fifo_level1 = (uart_rx_fifo_level0 + uart_rx_fifo_readable);
always @(*) begin
	uart_rx_fifo_wrport_adr = 4'd0;
	if (uart_rx_fifo_replace) begin
		uart_rx_fifo_wrport_adr = (uart_rx_fifo_produce - 1'd1);
	end else begin
		uart_rx_fifo_wrport_adr = uart_rx_fifo_produce;
	end
end
assign uart_rx_fifo_wrport_dat_w = uart_rx_fifo_syncfifo_din;
assign uart_rx_fifo_wrport_we = (uart_rx_fifo_syncfifo_we & (uart_rx_fifo_syncfifo_writable | uart_rx_fifo_replace));
assign uart_rx_fifo_do_read = (uart_rx_fifo_syncfifo_readable & uart_rx_fifo_syncfifo_re);
assign uart_rx_fifo_rdport_adr = uart_rx_fifo_consume;
assign uart_rx_fifo_syncfifo_dout = uart_rx_fifo_rdport_dat_r;
assign uart_rx_fifo_rdport_re = uart_rx_fifo_do_read;
assign uart_rx_fifo_syncfifo_writable = (uart_rx_fifo_level0 != 5'd16);
assign uart_rx_fifo_syncfifo_readable = (uart_rx_fifo_level0 != 1'd0);
assign dbg_uart_wait = (~dbg_uart_is_ongoing);
assign dbg_uart_reset = dbg_uart_done;
assign dbg_uart_wishbone_adr = dbg_uart_address;
assign dbg_uart_wishbone_dat_w = dbg_uart_data;
assign dbg_uart_wishbone_sel = 4'd15;
always @(*) begin
	dbg_uart_tx_sink_payload_data = 8'd0;
	case (dbg_uart_bytes_count)
		1'd0: begin
			dbg_uart_tx_sink_payload_data = dbg_uart_data[31:24];
		end
		1'd1: begin
			dbg_uart_tx_sink_payload_data = dbg_uart_data[31:16];
		end
		2'd2: begin
			dbg_uart_tx_sink_payload_data = dbg_uart_data[31:8];
		end
		2'd3: begin
			dbg_uart_tx_sink_payload_data = dbg_uart_data[31:0];
		end
	endcase
end
assign dbg_uart_tx_sink_last = ((dbg_uart_bytes_count == 2'd3) & (dbg_uart_words_count == (dbg_uart_length - 1'd1)));
always @(*) begin
	uartwishbonebridge_rs232phytx_next_state = 1'd0;
	uartwishbonebridge_rs232phytx_next_state = uartwishbonebridge_rs232phytx_state;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				if ((dbg_uart_tx_count == 4'd9)) begin
					uartwishbonebridge_rs232phytx_next_state = 1'd0;
				end
			end
		end
		default: begin
			if (dbg_uart_tx_sink_valid) begin
				uartwishbonebridge_rs232phytx_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_sink_ready = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				if ((dbg_uart_tx_count == 4'd9)) begin
					dbg_uart_tx_sink_ready = 1'd1;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2 = 8'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2 = {1'd1, dbg_uart_tx_data[7:1]};
			end
		end
		default: begin
			if (dbg_uart_tx_sink_valid) begin
				dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2 = dbg_uart_tx_sink_payload_data;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2 = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2 = 1'd1;
			end
		end
		default: begin
			if (dbg_uart_tx_sink_valid) begin
				dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_enable = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			dbg_uart_tx_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0 = 4'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0 = (dbg_uart_tx_count + 1'd1);
			end
		end
		default: begin
			dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0 = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = dbg_uart_tx_data;
			end
		end
		default: begin
			dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = 1'd1;
			if (dbg_uart_tx_sink_valid) begin
				dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1 = 1'd0;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd0;
	case (uartwishbonebridge_rs232phytx_state)
		1'd1: begin
			if (dbg_uart_tx_tick) begin
				dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd1;
			end
		end
		default: begin
			dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd1;
			if (dbg_uart_tx_sink_valid) begin
				dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	uartwishbonebridge_rs232phyrx_next_state = 1'd0;
	uartwishbonebridge_rs232phyrx_next_state = uartwishbonebridge_rs232phyrx_state;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				if ((dbg_uart_rx_count == 4'd9)) begin
					uartwishbonebridge_rs232phyrx_next_state = 1'd0;
				end
			end
		end
		default: begin
			if (((dbg_uart_rx_rx == 1'd0) & (dbg_uart_rx_rx_d == 1'd1))) begin
				uartwishbonebridge_rs232phyrx_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_source_valid = 1'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				if ((dbg_uart_rx_count == 4'd9)) begin
					dbg_uart_rx_source_valid = (dbg_uart_rx_rx == 1'd1);
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value1 = 8'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value1 = {dbg_uart_rx_rx, dbg_uart_rx_data[7:1]};
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value_ce1 = 1'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value_ce1 = 1'd1;
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_source_payload_data = 8'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				if ((dbg_uart_rx_count == 4'd9)) begin
					dbg_uart_rx_source_payload_data = dbg_uart_rx_data;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_enable = 1'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			dbg_uart_rx_enable = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0 = 4'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0 = (dbg_uart_rx_count + 1'd1);
			end
		end
		default: begin
			dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0 = 1'd0;
	case (uartwishbonebridge_rs232phyrx_state)
		1'd1: begin
			if (dbg_uart_rx_tick) begin
				dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	uartwishbonebridge_next_state = 3'd0;
	uartwishbonebridge_next_state = uartwishbonebridge_state;
	case (uartwishbonebridge_state)
		1'd1: begin
			if (dbg_uart_rx_source_valid) begin
				uartwishbonebridge_next_state = 2'd2;
			end
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					if (((dbg_uart_cmd == 1'd1) | (dbg_uart_cmd == 2'd3))) begin
						uartwishbonebridge_next_state = 2'd3;
					end else begin
						if (((dbg_uart_cmd == 2'd2) | (dbg_uart_cmd == 3'd4))) begin
							uartwishbonebridge_next_state = 3'd5;
						end else begin
							uartwishbonebridge_next_state = 1'd0;
						end
					end
				end
			end
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					uartwishbonebridge_next_state = 3'd4;
				end
			end
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				if ((dbg_uart_words_count == (dbg_uart_length - 1'd1))) begin
					uartwishbonebridge_next_state = 1'd0;
				end else begin
					uartwishbonebridge_next_state = 2'd3;
				end
			end
		end
		3'd5: begin
			if (dbg_uart_wishbone_ack) begin
				uartwishbonebridge_next_state = 3'd6;
			end
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					if ((dbg_uart_words_count == (dbg_uart_length - 1'd1))) begin
						uartwishbonebridge_next_state = 1'd0;
					end else begin
						uartwishbonebridge_next_state = 3'd5;
					end
				end
			end
		end
		default: begin
			if (dbg_uart_rx_source_valid) begin
				uartwishbonebridge_next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_bytes_count_uartwishbonebridge_next_value0 = 2'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value0 = (dbg_uart_bytes_count + 1'd1);
			end
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value0 = (dbg_uart_bytes_count + 1'd1);
			end
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value0 = (dbg_uart_bytes_count + 1'd1);
			end
		end
		default: begin
			dbg_uart_bytes_count_uartwishbonebridge_next_value0 = 1'd0;
		end
	endcase
end
always @(*) begin
	dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd1;
			end
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd1;
			end
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd1;
			end
		end
		default: begin
			dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0 = 1'd1;
		end
	endcase
end
always @(*) begin
	dbg_uart_wishbone_cyc = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			dbg_uart_wishbone_cyc = 1'd1;
		end
		3'd5: begin
			dbg_uart_wishbone_cyc = 1'd1;
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_wishbone_stb = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			dbg_uart_wishbone_stb = 1'd1;
		end
		3'd5: begin
			dbg_uart_wishbone_stb = 1'd1;
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_words_count_uartwishbonebridge_next_value1 = 8'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_words_count_uartwishbonebridge_next_value1 = (dbg_uart_words_count + 1'd1);
			end
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					dbg_uart_words_count_uartwishbonebridge_next_value1 = (dbg_uart_words_count + 1'd1);
				end
			end
		end
		default: begin
			dbg_uart_words_count_uartwishbonebridge_next_value1 = 1'd0;
		end
	endcase
end
always @(*) begin
	dbg_uart_wishbone_we = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			dbg_uart_wishbone_we = 1'd1;
		end
		3'd5: begin
			dbg_uart_wishbone_we = 1'd0;
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd1;
			end
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd1;
				end
			end
		end
		default: begin
			dbg_uart_words_count_uartwishbonebridge_next_value_ce1 = 1'd1;
		end
	endcase
end
always @(*) begin
	dbg_uart_cmd_uartwishbonebridge_next_value2 = 8'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_cmd_uartwishbonebridge_next_value2 = dbg_uart_rx_source_payload_data;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_cmd_uartwishbonebridge_next_value_ce2 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_cmd_uartwishbonebridge_next_value_ce2 = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	dbg_uart_length_uartwishbonebridge_next_value3 = 8'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_length_uartwishbonebridge_next_value3 = dbg_uart_rx_source_payload_data;
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_length_uartwishbonebridge_next_value_ce3 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_length_uartwishbonebridge_next_value_ce3 = 1'd1;
			end
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_address_uartwishbonebridge_next_value4 = 32'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_address_uartwishbonebridge_next_value4 = {dbg_uart_address, dbg_uart_rx_source_payload_data};
			end
		end
		2'd3: begin
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_address_uartwishbonebridge_next_value4 = (dbg_uart_address + dbg_uart_incr);
			end
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					dbg_uart_address_uartwishbonebridge_next_value4 = (dbg_uart_address + dbg_uart_incr);
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd1;
			end
		end
		2'd3: begin
		end
		3'd4: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd1;
			end
		end
		3'd5: begin
		end
		3'd6: begin
			if (dbg_uart_tx_sink_ready) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					dbg_uart_address_uartwishbonebridge_next_value_ce4 = 1'd1;
				end
			end
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_incr_uartwishbonebridge_next_value5 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					if (((dbg_uart_cmd == 1'd1) | (dbg_uart_cmd == 2'd3))) begin
						dbg_uart_incr_uartwishbonebridge_next_value5 = (dbg_uart_cmd == 1'd1);
					end else begin
						if (((dbg_uart_cmd == 2'd2) | (dbg_uart_cmd == 3'd4))) begin
							dbg_uart_incr_uartwishbonebridge_next_value5 = (dbg_uart_cmd == 2'd2);
						end else begin
						end
					end
				end
			end
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_incr_uartwishbonebridge_next_value_ce5 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
			if (dbg_uart_rx_source_valid) begin
				if ((dbg_uart_bytes_count == 2'd3)) begin
					if (((dbg_uart_cmd == 1'd1) | (dbg_uart_cmd == 2'd3))) begin
						dbg_uart_incr_uartwishbonebridge_next_value_ce5 = 1'd1;
					end else begin
						if (((dbg_uart_cmd == 2'd2) | (dbg_uart_cmd == 3'd4))) begin
							dbg_uart_incr_uartwishbonebridge_next_value_ce5 = 1'd1;
						end else begin
						end
					end
				end
			end
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_tx_sink_valid = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
			dbg_uart_tx_sink_valid = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_data_uartwishbonebridge_next_value6 = 32'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_data_uartwishbonebridge_next_value6 = {dbg_uart_data, dbg_uart_rx_source_payload_data};
			end
		end
		3'd4: begin
		end
		3'd5: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_data_uartwishbonebridge_next_value6 = dbg_uart_wishbone_dat_r;
			end
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_is_ongoing = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
		end
		3'd4: begin
		end
		3'd5: begin
		end
		3'd6: begin
		end
		default: begin
			dbg_uart_is_ongoing = 1'd1;
		end
	endcase
end
always @(*) begin
	dbg_uart_data_uartwishbonebridge_next_value_ce6 = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
		end
		2'd2: begin
		end
		2'd3: begin
			if (dbg_uart_rx_source_valid) begin
				dbg_uart_data_uartwishbonebridge_next_value_ce6 = 1'd1;
			end
		end
		3'd4: begin
		end
		3'd5: begin
			if (dbg_uart_wishbone_ack) begin
				dbg_uart_data_uartwishbonebridge_next_value_ce6 = 1'd1;
			end
		end
		3'd6: begin
		end
		default: begin
		end
	endcase
end
always @(*) begin
	dbg_uart_rx_source_ready = 1'd0;
	case (uartwishbonebridge_state)
		1'd1: begin
			dbg_uart_rx_source_ready = 1'd1;
		end
		2'd2: begin
			dbg_uart_rx_source_ready = 1'd1;
		end
		2'd3: begin
			dbg_uart_rx_source_ready = 1'd1;
		end
		3'd4: begin
			dbg_uart_rx_source_ready = 1'd0;
		end
		3'd5: begin
			dbg_uart_rx_source_ready = 1'd0;
		end
		3'd6: begin
			dbg_uart_rx_source_ready = 1'd0;
		end
		default: begin
			dbg_uart_rx_source_ready = 1'd1;
		end
	endcase
end
assign dbg_uart_done = (dbg_uart_count == 1'd0);
assign debug_oeb = debug_oeb_storage;
assign debug_mode = debug_mode_storage;
assign uart_enabled_o = uart_enabled_storage;
assign gpio_mode0_pad = gpio_mode0_storage;
assign gpio_mode1_pad = gpio_mode1_storage;
assign gpio_inenb_pad = (~gpio_ien_storage);
assign gpio_outenb_pad = (~gpio_oe_storage);
assign gpio_out_pad = gpio_out_storage;
always @(*) begin
	la_iena = 128'd0;
	la_iena[0] = (~la_ien_storage[0]);
	la_iena[1] = (~la_ien_storage[1]);
	la_iena[2] = (~la_ien_storage[2]);
	la_iena[3] = (~la_ien_storage[3]);
	la_iena[4] = (~la_ien_storage[4]);
	la_iena[5] = (~la_ien_storage[5]);
	la_iena[6] = (~la_ien_storage[6]);
	la_iena[7] = (~la_ien_storage[7]);
	la_iena[8] = (~la_ien_storage[8]);
	la_iena[9] = (~la_ien_storage[9]);
	la_iena[10] = (~la_ien_storage[10]);
	la_iena[11] = (~la_ien_storage[11]);
	la_iena[12] = (~la_ien_storage[12]);
	la_iena[13] = (~la_ien_storage[13]);
	la_iena[14] = (~la_ien_storage[14]);
	la_iena[15] = (~la_ien_storage[15]);
	la_iena[16] = (~la_ien_storage[16]);
	la_iena[17] = (~la_ien_storage[17]);
	la_iena[18] = (~la_ien_storage[18]);
	la_iena[19] = (~la_ien_storage[19]);
	la_iena[20] = (~la_ien_storage[20]);
	la_iena[21] = (~la_ien_storage[21]);
	la_iena[22] = (~la_ien_storage[22]);
	la_iena[23] = (~la_ien_storage[23]);
	la_iena[24] = (~la_ien_storage[24]);
	la_iena[25] = (~la_ien_storage[25]);
	la_iena[26] = (~la_ien_storage[26]);
	la_iena[27] = (~la_ien_storage[27]);
	la_iena[28] = (~la_ien_storage[28]);
	la_iena[29] = (~la_ien_storage[29]);
	la_iena[30] = (~la_ien_storage[30]);
	la_iena[31] = (~la_ien_storage[31]);
	la_iena[32] = (~la_ien_storage[32]);
	la_iena[33] = (~la_ien_storage[33]);
	la_iena[34] = (~la_ien_storage[34]);
	la_iena[35] = (~la_ien_storage[35]);
	la_iena[36] = (~la_ien_storage[36]);
	la_iena[37] = (~la_ien_storage[37]);
	la_iena[38] = (~la_ien_storage[38]);
	la_iena[39] = (~la_ien_storage[39]);
	la_iena[40] = (~la_ien_storage[40]);
	la_iena[41] = (~la_ien_storage[41]);
	la_iena[42] = (~la_ien_storage[42]);
	la_iena[43] = (~la_ien_storage[43]);
	la_iena[44] = (~la_ien_storage[44]);
	la_iena[45] = (~la_ien_storage[45]);
	la_iena[46] = (~la_ien_storage[46]);
	la_iena[47] = (~la_ien_storage[47]);
	la_iena[48] = (~la_ien_storage[48]);
	la_iena[49] = (~la_ien_storage[49]);
	la_iena[50] = (~la_ien_storage[50]);
	la_iena[51] = (~la_ien_storage[51]);
	la_iena[52] = (~la_ien_storage[52]);
	la_iena[53] = (~la_ien_storage[53]);
	la_iena[54] = (~la_ien_storage[54]);
	la_iena[55] = (~la_ien_storage[55]);
	la_iena[56] = (~la_ien_storage[56]);
	la_iena[57] = (~la_ien_storage[57]);
	la_iena[58] = (~la_ien_storage[58]);
	la_iena[59] = (~la_ien_storage[59]);
	la_iena[60] = (~la_ien_storage[60]);
	la_iena[61] = (~la_ien_storage[61]);
	la_iena[62] = (~la_ien_storage[62]);
	la_iena[63] = (~la_ien_storage[63]);
	la_iena[64] = (~la_ien_storage[64]);
	la_iena[65] = (~la_ien_storage[65]);
	la_iena[66] = (~la_ien_storage[66]);
	la_iena[67] = (~la_ien_storage[67]);
	la_iena[68] = (~la_ien_storage[68]);
	la_iena[69] = (~la_ien_storage[69]);
	la_iena[70] = (~la_ien_storage[70]);
	la_iena[71] = (~la_ien_storage[71]);
	la_iena[72] = (~la_ien_storage[72]);
	la_iena[73] = (~la_ien_storage[73]);
	la_iena[74] = (~la_ien_storage[74]);
	la_iena[75] = (~la_ien_storage[75]);
	la_iena[76] = (~la_ien_storage[76]);
	la_iena[77] = (~la_ien_storage[77]);
	la_iena[78] = (~la_ien_storage[78]);
	la_iena[79] = (~la_ien_storage[79]);
	la_iena[80] = (~la_ien_storage[80]);
	la_iena[81] = (~la_ien_storage[81]);
	la_iena[82] = (~la_ien_storage[82]);
	la_iena[83] = (~la_ien_storage[83]);
	la_iena[84] = (~la_ien_storage[84]);
	la_iena[85] = (~la_ien_storage[85]);
	la_iena[86] = (~la_ien_storage[86]);
	la_iena[87] = (~la_ien_storage[87]);
	la_iena[88] = (~la_ien_storage[88]);
	la_iena[89] = (~la_ien_storage[89]);
	la_iena[90] = (~la_ien_storage[90]);
	la_iena[91] = (~la_ien_storage[91]);
	la_iena[92] = (~la_ien_storage[92]);
	la_iena[93] = (~la_ien_storage[93]);
	la_iena[94] = (~la_ien_storage[94]);
	la_iena[95] = (~la_ien_storage[95]);
	la_iena[96] = (~la_ien_storage[96]);
	la_iena[97] = (~la_ien_storage[97]);
	la_iena[98] = (~la_ien_storage[98]);
	la_iena[99] = (~la_ien_storage[99]);
	la_iena[100] = (~la_ien_storage[100]);
	la_iena[101] = (~la_ien_storage[101]);
	la_iena[102] = (~la_ien_storage[102]);
	la_iena[103] = (~la_ien_storage[103]);
	la_iena[104] = (~la_ien_storage[104]);
	la_iena[105] = (~la_ien_storage[105]);
	la_iena[106] = (~la_ien_storage[106]);
	la_iena[107] = (~la_ien_storage[107]);
	la_iena[108] = (~la_ien_storage[108]);
	la_iena[109] = (~la_ien_storage[109]);
	la_iena[110] = (~la_ien_storage[110]);
	la_iena[111] = (~la_ien_storage[111]);
	la_iena[112] = (~la_ien_storage[112]);
	la_iena[113] = (~la_ien_storage[113]);
	la_iena[114] = (~la_ien_storage[114]);
	la_iena[115] = (~la_ien_storage[115]);
	la_iena[116] = (~la_ien_storage[116]);
	la_iena[117] = (~la_ien_storage[117]);
	la_iena[118] = (~la_ien_storage[118]);
	la_iena[119] = (~la_ien_storage[119]);
	la_iena[120] = (~la_ien_storage[120]);
	la_iena[121] = (~la_ien_storage[121]);
	la_iena[122] = (~la_ien_storage[122]);
	la_iena[123] = (~la_ien_storage[123]);
	la_iena[124] = (~la_ien_storage[124]);
	la_iena[125] = (~la_ien_storage[125]);
	la_iena[126] = (~la_ien_storage[126]);
	la_iena[127] = (~la_ien_storage[127]);
end
always @(*) begin
	la_oenb = 128'd0;
	la_oenb[0] = (~la_oe_storage[0]);
	la_oenb[1] = (~la_oe_storage[1]);
	la_oenb[2] = (~la_oe_storage[2]);
	la_oenb[3] = (~la_oe_storage[3]);
	la_oenb[4] = (~la_oe_storage[4]);
	la_oenb[5] = (~la_oe_storage[5]);
	la_oenb[6] = (~la_oe_storage[6]);
	la_oenb[7] = (~la_oe_storage[7]);
	la_oenb[8] = (~la_oe_storage[8]);
	la_oenb[9] = (~la_oe_storage[9]);
	la_oenb[10] = (~la_oe_storage[10]);
	la_oenb[11] = (~la_oe_storage[11]);
	la_oenb[12] = (~la_oe_storage[12]);
	la_oenb[13] = (~la_oe_storage[13]);
	la_oenb[14] = (~la_oe_storage[14]);
	la_oenb[15] = (~la_oe_storage[15]);
	la_oenb[16] = (~la_oe_storage[16]);
	la_oenb[17] = (~la_oe_storage[17]);
	la_oenb[18] = (~la_oe_storage[18]);
	la_oenb[19] = (~la_oe_storage[19]);
	la_oenb[20] = (~la_oe_storage[20]);
	la_oenb[21] = (~la_oe_storage[21]);
	la_oenb[22] = (~la_oe_storage[22]);
	la_oenb[23] = (~la_oe_storage[23]);
	la_oenb[24] = (~la_oe_storage[24]);
	la_oenb[25] = (~la_oe_storage[25]);
	la_oenb[26] = (~la_oe_storage[26]);
	la_oenb[27] = (~la_oe_storage[27]);
	la_oenb[28] = (~la_oe_storage[28]);
	la_oenb[29] = (~la_oe_storage[29]);
	la_oenb[30] = (~la_oe_storage[30]);
	la_oenb[31] = (~la_oe_storage[31]);
	la_oenb[32] = (~la_oe_storage[32]);
	la_oenb[33] = (~la_oe_storage[33]);
	la_oenb[34] = (~la_oe_storage[34]);
	la_oenb[35] = (~la_oe_storage[35]);
	la_oenb[36] = (~la_oe_storage[36]);
	la_oenb[37] = (~la_oe_storage[37]);
	la_oenb[38] = (~la_oe_storage[38]);
	la_oenb[39] = (~la_oe_storage[39]);
	la_oenb[40] = (~la_oe_storage[40]);
	la_oenb[41] = (~la_oe_storage[41]);
	la_oenb[42] = (~la_oe_storage[42]);
	la_oenb[43] = (~la_oe_storage[43]);
	la_oenb[44] = (~la_oe_storage[44]);
	la_oenb[45] = (~la_oe_storage[45]);
	la_oenb[46] = (~la_oe_storage[46]);
	la_oenb[47] = (~la_oe_storage[47]);
	la_oenb[48] = (~la_oe_storage[48]);
	la_oenb[49] = (~la_oe_storage[49]);
	la_oenb[50] = (~la_oe_storage[50]);
	la_oenb[51] = (~la_oe_storage[51]);
	la_oenb[52] = (~la_oe_storage[52]);
	la_oenb[53] = (~la_oe_storage[53]);
	la_oenb[54] = (~la_oe_storage[54]);
	la_oenb[55] = (~la_oe_storage[55]);
	la_oenb[56] = (~la_oe_storage[56]);
	la_oenb[57] = (~la_oe_storage[57]);
	la_oenb[58] = (~la_oe_storage[58]);
	la_oenb[59] = (~la_oe_storage[59]);
	la_oenb[60] = (~la_oe_storage[60]);
	la_oenb[61] = (~la_oe_storage[61]);
	la_oenb[62] = (~la_oe_storage[62]);
	la_oenb[63] = (~la_oe_storage[63]);
	la_oenb[64] = (~la_oe_storage[64]);
	la_oenb[65] = (~la_oe_storage[65]);
	la_oenb[66] = (~la_oe_storage[66]);
	la_oenb[67] = (~la_oe_storage[67]);
	la_oenb[68] = (~la_oe_storage[68]);
	la_oenb[69] = (~la_oe_storage[69]);
	la_oenb[70] = (~la_oe_storage[70]);
	la_oenb[71] = (~la_oe_storage[71]);
	la_oenb[72] = (~la_oe_storage[72]);
	la_oenb[73] = (~la_oe_storage[73]);
	la_oenb[74] = (~la_oe_storage[74]);
	la_oenb[75] = (~la_oe_storage[75]);
	la_oenb[76] = (~la_oe_storage[76]);
	la_oenb[77] = (~la_oe_storage[77]);
	la_oenb[78] = (~la_oe_storage[78]);
	la_oenb[79] = (~la_oe_storage[79]);
	la_oenb[80] = (~la_oe_storage[80]);
	la_oenb[81] = (~la_oe_storage[81]);
	la_oenb[82] = (~la_oe_storage[82]);
	la_oenb[83] = (~la_oe_storage[83]);
	la_oenb[84] = (~la_oe_storage[84]);
	la_oenb[85] = (~la_oe_storage[85]);
	la_oenb[86] = (~la_oe_storage[86]);
	la_oenb[87] = (~la_oe_storage[87]);
	la_oenb[88] = (~la_oe_storage[88]);
	la_oenb[89] = (~la_oe_storage[89]);
	la_oenb[90] = (~la_oe_storage[90]);
	la_oenb[91] = (~la_oe_storage[91]);
	la_oenb[92] = (~la_oe_storage[92]);
	la_oenb[93] = (~la_oe_storage[93]);
	la_oenb[94] = (~la_oe_storage[94]);
	la_oenb[95] = (~la_oe_storage[95]);
	la_oenb[96] = (~la_oe_storage[96]);
	la_oenb[97] = (~la_oe_storage[97]);
	la_oenb[98] = (~la_oe_storage[98]);
	la_oenb[99] = (~la_oe_storage[99]);
	la_oenb[100] = (~la_oe_storage[100]);
	la_oenb[101] = (~la_oe_storage[101]);
	la_oenb[102] = (~la_oe_storage[102]);
	la_oenb[103] = (~la_oe_storage[103]);
	la_oenb[104] = (~la_oe_storage[104]);
	la_oenb[105] = (~la_oe_storage[105]);
	la_oenb[106] = (~la_oe_storage[106]);
	la_oenb[107] = (~la_oe_storage[107]);
	la_oenb[108] = (~la_oe_storage[108]);
	la_oenb[109] = (~la_oe_storage[109]);
	la_oenb[110] = (~la_oe_storage[110]);
	la_oenb[111] = (~la_oe_storage[111]);
	la_oenb[112] = (~la_oe_storage[112]);
	la_oenb[113] = (~la_oe_storage[113]);
	la_oenb[114] = (~la_oe_storage[114]);
	la_oenb[115] = (~la_oe_storage[115]);
	la_oenb[116] = (~la_oe_storage[116]);
	la_oenb[117] = (~la_oe_storage[117]);
	la_oenb[118] = (~la_oe_storage[118]);
	la_oenb[119] = (~la_oe_storage[119]);
	la_oenb[120] = (~la_oe_storage[120]);
	la_oenb[121] = (~la_oe_storage[121]);
	la_oenb[122] = (~la_oe_storage[122]);
	la_oenb[123] = (~la_oe_storage[123]);
	la_oenb[124] = (~la_oe_storage[124]);
	la_oenb[125] = (~la_oe_storage[125]);
	la_oenb[126] = (~la_oe_storage[126]);
	la_oenb[127] = (~la_oe_storage[127]);
end
always @(*) begin
	la_output = 128'd0;
	la_output[0] = la_out_storage[0];
	la_output[1] = la_out_storage[1];
	la_output[2] = la_out_storage[2];
	la_output[3] = la_out_storage[3];
	la_output[4] = la_out_storage[4];
	la_output[5] = la_out_storage[5];
	la_output[6] = la_out_storage[6];
	la_output[7] = la_out_storage[7];
	la_output[8] = la_out_storage[8];
	la_output[9] = la_out_storage[9];
	la_output[10] = la_out_storage[10];
	la_output[11] = la_out_storage[11];
	la_output[12] = la_out_storage[12];
	la_output[13] = la_out_storage[13];
	la_output[14] = la_out_storage[14];
	la_output[15] = la_out_storage[15];
	la_output[16] = la_out_storage[16];
	la_output[17] = la_out_storage[17];
	la_output[18] = la_out_storage[18];
	la_output[19] = la_out_storage[19];
	la_output[20] = la_out_storage[20];
	la_output[21] = la_out_storage[21];
	la_output[22] = la_out_storage[22];
	la_output[23] = la_out_storage[23];
	la_output[24] = la_out_storage[24];
	la_output[25] = la_out_storage[25];
	la_output[26] = la_out_storage[26];
	la_output[27] = la_out_storage[27];
	la_output[28] = la_out_storage[28];
	la_output[29] = la_out_storage[29];
	la_output[30] = la_out_storage[30];
	la_output[31] = la_out_storage[31];
	la_output[32] = la_out_storage[32];
	la_output[33] = la_out_storage[33];
	la_output[34] = la_out_storage[34];
	la_output[35] = la_out_storage[35];
	la_output[36] = la_out_storage[36];
	la_output[37] = la_out_storage[37];
	la_output[38] = la_out_storage[38];
	la_output[39] = la_out_storage[39];
	la_output[40] = la_out_storage[40];
	la_output[41] = la_out_storage[41];
	la_output[42] = la_out_storage[42];
	la_output[43] = la_out_storage[43];
	la_output[44] = la_out_storage[44];
	la_output[45] = la_out_storage[45];
	la_output[46] = la_out_storage[46];
	la_output[47] = la_out_storage[47];
	la_output[48] = la_out_storage[48];
	la_output[49] = la_out_storage[49];
	la_output[50] = la_out_storage[50];
	la_output[51] = la_out_storage[51];
	la_output[52] = la_out_storage[52];
	la_output[53] = la_out_storage[53];
	la_output[54] = la_out_storage[54];
	la_output[55] = la_out_storage[55];
	la_output[56] = la_out_storage[56];
	la_output[57] = la_out_storage[57];
	la_output[58] = la_out_storage[58];
	la_output[59] = la_out_storage[59];
	la_output[60] = la_out_storage[60];
	la_output[61] = la_out_storage[61];
	la_output[62] = la_out_storage[62];
	la_output[63] = la_out_storage[63];
	la_output[64] = la_out_storage[64];
	la_output[65] = la_out_storage[65];
	la_output[66] = la_out_storage[66];
	la_output[67] = la_out_storage[67];
	la_output[68] = la_out_storage[68];
	la_output[69] = la_out_storage[69];
	la_output[70] = la_out_storage[70];
	la_output[71] = la_out_storage[71];
	la_output[72] = la_out_storage[72];
	la_output[73] = la_out_storage[73];
	la_output[74] = la_out_storage[74];
	la_output[75] = la_out_storage[75];
	la_output[76] = la_out_storage[76];
	la_output[77] = la_out_storage[77];
	la_output[78] = la_out_storage[78];
	la_output[79] = la_out_storage[79];
	la_output[80] = la_out_storage[80];
	la_output[81] = la_out_storage[81];
	la_output[82] = la_out_storage[82];
	la_output[83] = la_out_storage[83];
	la_output[84] = la_out_storage[84];
	la_output[85] = la_out_storage[85];
	la_output[86] = la_out_storage[86];
	la_output[87] = la_out_storage[87];
	la_output[88] = la_out_storage[88];
	la_output[89] = la_out_storage[89];
	la_output[90] = la_out_storage[90];
	la_output[91] = la_out_storage[91];
	la_output[92] = la_out_storage[92];
	la_output[93] = la_out_storage[93];
	la_output[94] = la_out_storage[94];
	la_output[95] = la_out_storage[95];
	la_output[96] = la_out_storage[96];
	la_output[97] = la_out_storage[97];
	la_output[98] = la_out_storage[98];
	la_output[99] = la_out_storage[99];
	la_output[100] = la_out_storage[100];
	la_output[101] = la_out_storage[101];
	la_output[102] = la_out_storage[102];
	la_output[103] = la_out_storage[103];
	la_output[104] = la_out_storage[104];
	la_output[105] = la_out_storage[105];
	la_output[106] = la_out_storage[106];
	la_output[107] = la_out_storage[107];
	la_output[108] = la_out_storage[108];
	la_output[109] = la_out_storage[109];
	la_output[110] = la_out_storage[110];
	la_output[111] = la_out_storage[111];
	la_output[112] = la_out_storage[112];
	la_output[113] = la_out_storage[113];
	la_output[114] = la_out_storage[114];
	la_output[115] = la_out_storage[115];
	la_output[116] = la_out_storage[116];
	la_output[117] = la_out_storage[117];
	la_output[118] = la_out_storage[118];
	la_output[119] = la_out_storage[119];
	la_output[120] = la_out_storage[120];
	la_output[121] = la_out_storage[121];
	la_output[122] = la_out_storage[122];
	la_output[123] = la_out_storage[123];
	la_output[124] = la_out_storage[124];
	la_output[125] = la_out_storage[125];
	la_output[126] = la_out_storage[126];
	la_output[127] = la_out_storage[127];
end
assign spi_enabled = spi_enabled_storage;
assign user_irq_ena = user_irq_ena_storage;
always @(*) begin
	gpioin0_gpioin0_trigger = 1'd0;
	if (gpioin0_gpioin0_mode_storage) begin
		gpioin0_gpioin0_trigger = (gpioin0_in_status ^ gpioin0_gpioin0_in_pads_n_d);
	end else begin
		gpioin0_gpioin0_trigger = (gpioin0_in_status ^ gpioin0_gpioin0_edge_storage);
	end
end
assign gpioin0_i00 = gpioin0_gpioin0_status;
assign gpioin0_i01 = gpioin0_gpioin0_pending;
always @(*) begin
	gpioin0_gpioin0_clear = 1'd0;
	if ((gpioin0_pending_re & gpioin0_pending_r)) begin
		gpioin0_gpioin0_clear = 1'd1;
	end
end
assign gpioin0_gpioin0_irq = (gpioin0_pending_status & gpioin0_enable_storage);
assign gpioin0_gpioin0_status = gpioin0_gpioin0_trigger;
always @(*) begin
	gpioin1_gpioin1_trigger = 1'd0;
	if (gpioin1_gpioin1_mode_storage) begin
		gpioin1_gpioin1_trigger = (gpioin1_in_status ^ gpioin1_gpioin1_in_pads_n_d);
	end else begin
		gpioin1_gpioin1_trigger = (gpioin1_in_status ^ gpioin1_gpioin1_edge_storage);
	end
end
assign gpioin1_i00 = gpioin1_gpioin1_status;
assign gpioin1_i01 = gpioin1_gpioin1_pending;
always @(*) begin
	gpioin1_gpioin1_clear = 1'd0;
	if ((gpioin1_pending_re & gpioin1_pending_r)) begin
		gpioin1_gpioin1_clear = 1'd1;
	end
end
assign gpioin1_gpioin1_irq = (gpioin1_pending_status & gpioin1_enable_storage);
assign gpioin1_gpioin1_status = gpioin1_gpioin1_trigger;
always @(*) begin
	gpioin2_gpioin2_trigger = 1'd0;
	if (gpioin2_gpioin2_mode_storage) begin
		gpioin2_gpioin2_trigger = (gpioin2_in_status ^ gpioin2_gpioin2_in_pads_n_d);
	end else begin
		gpioin2_gpioin2_trigger = (gpioin2_in_status ^ gpioin2_gpioin2_edge_storage);
	end
end
assign gpioin2_i00 = gpioin2_gpioin2_status;
assign gpioin2_i01 = gpioin2_gpioin2_pending;
always @(*) begin
	gpioin2_gpioin2_clear = 1'd0;
	if ((gpioin2_pending_re & gpioin2_pending_r)) begin
		gpioin2_gpioin2_clear = 1'd1;
	end
end
assign gpioin2_gpioin2_irq = (gpioin2_pending_status & gpioin2_enable_storage);
assign gpioin2_gpioin2_status = gpioin2_gpioin2_trigger;
always @(*) begin
	gpioin3_gpioin3_trigger = 1'd0;
	if (gpioin3_gpioin3_mode_storage) begin
		gpioin3_gpioin3_trigger = (gpioin3_in_status ^ gpioin3_gpioin3_in_pads_n_d);
	end else begin
		gpioin3_gpioin3_trigger = (gpioin3_in_status ^ gpioin3_gpioin3_edge_storage);
	end
end
assign gpioin3_i00 = gpioin3_gpioin3_status;
assign gpioin3_i01 = gpioin3_gpioin3_pending;
always @(*) begin
	gpioin3_gpioin3_clear = 1'd0;
	if ((gpioin3_pending_re & gpioin3_pending_r)) begin
		gpioin3_gpioin3_clear = 1'd1;
	end
end
assign gpioin3_gpioin3_irq = (gpioin3_pending_status & gpioin3_enable_storage);
assign gpioin3_gpioin3_status = gpioin3_gpioin3_trigger;
always @(*) begin
	gpioin4_gpioin4_trigger = 1'd0;
	if (gpioin4_gpioin4_mode_storage) begin
		gpioin4_gpioin4_trigger = (gpioin4_in_status ^ gpioin4_gpioin4_in_pads_n_d);
	end else begin
		gpioin4_gpioin4_trigger = (gpioin4_in_status ^ gpioin4_gpioin4_edge_storage);
	end
end
assign gpioin4_i00 = gpioin4_gpioin4_status;
assign gpioin4_i01 = gpioin4_gpioin4_pending;
always @(*) begin
	gpioin4_gpioin4_clear = 1'd0;
	if ((gpioin4_pending_re & gpioin4_pending_r)) begin
		gpioin4_gpioin4_clear = 1'd1;
	end
end
assign gpioin4_gpioin4_irq = (gpioin4_pending_status & gpioin4_enable_storage);
assign gpioin4_gpioin4_status = gpioin4_gpioin4_trigger;
always @(*) begin
	gpioin5_gpioin5_trigger = 1'd0;
	if (gpioin5_gpioin5_mode_storage) begin
		gpioin5_gpioin5_trigger = (gpioin5_in_status ^ gpioin5_gpioin5_in_pads_n_d);
	end else begin
		gpioin5_gpioin5_trigger = (gpioin5_in_status ^ gpioin5_gpioin5_edge_storage);
	end
end
assign gpioin5_i00 = gpioin5_gpioin5_status;
assign gpioin5_i01 = gpioin5_gpioin5_pending;
always @(*) begin
	gpioin5_gpioin5_clear = 1'd0;
	if ((gpioin5_pending_re & gpioin5_pending_r)) begin
		gpioin5_gpioin5_clear = 1'd1;
	end
end
assign gpioin5_gpioin5_irq = (gpioin5_pending_status & gpioin5_enable_storage);
assign gpioin5_gpioin5_status = gpioin5_gpioin5_trigger;
always @(*) begin
	next_state = 1'd0;
	next_state = state;
	case (state)
		1'd1: begin
			next_state = 1'd0;
		end
		default: begin
			if ((mgmtsoc_wishbone_cyc & mgmtsoc_wishbone_stb)) begin
				next_state = 1'd1;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_dat_w = 32'd0;
	case (state)
		1'd1: begin
		end
		default: begin
			mgmtsoc_dat_w = mgmtsoc_wishbone_dat_w;
		end
	endcase
end
always @(*) begin
	mgmtsoc_wishbone_dat_r = 32'd0;
	case (state)
		1'd1: begin
			mgmtsoc_wishbone_dat_r = mgmtsoc_dat_r;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_wishbone_ack = 1'd0;
	case (state)
		1'd1: begin
			mgmtsoc_wishbone_ack = 1'd1;
		end
		default: begin
		end
	endcase
end
always @(*) begin
	mgmtsoc_adr = 14'd0;
	case (state)
		1'd1: begin
		end
		default: begin
			if ((mgmtsoc_wishbone_cyc & mgmtsoc_wishbone_stb)) begin
				mgmtsoc_adr = mgmtsoc_wishbone_adr;
			end
		end
	endcase
end
always @(*) begin
	mgmtsoc_we = 1'd0;
	case (state)
		1'd1: begin
		end
		default: begin
			if ((mgmtsoc_wishbone_cyc & mgmtsoc_wishbone_stb)) begin
				mgmtsoc_we = (mgmtsoc_wishbone_we & (mgmtsoc_wishbone_sel != 1'd0));
			end
		end
	endcase
end
assign shared_adr = comb_array_muxed0;
assign shared_dat_w = comb_array_muxed1;
assign shared_sel = comb_array_muxed2;
assign shared_cyc = comb_array_muxed3;
assign shared_stb = comb_array_muxed4;
assign shared_we = comb_array_muxed5;
assign shared_cti = comb_array_muxed6;
assign shared_bte = comb_array_muxed7;
assign mgmtsoc_ibus_ibus_dat_r = shared_dat_r;
assign mgmtsoc_dbus_dbus_dat_r = shared_dat_r;
assign dbg_uart_wishbone_dat_r = shared_dat_r;
assign mgmtsoc_ibus_ibus_ack = (shared_ack & (grant == 1'd0));
assign mgmtsoc_dbus_dbus_ack = (shared_ack & (grant == 1'd1));
assign dbg_uart_wishbone_ack = (shared_ack & (grant == 2'd2));
assign mgmtsoc_ibus_ibus_err = (shared_err & (grant == 1'd0));
assign mgmtsoc_dbus_dbus_err = (shared_err & (grant == 1'd1));
assign dbg_uart_wishbone_err = (shared_err & (grant == 2'd2));
assign request = {dbg_uart_wishbone_cyc, mgmtsoc_dbus_dbus_cyc, mgmtsoc_ibus_ibus_cyc};
always @(*) begin
	slave_sel = 7'd0;
	slave_sel[0] = (shared_adr[29:6] == 24'd15732480);
	slave_sel[1] = (shared_adr[29:8] == 1'd0);
	slave_sel[2] = (shared_adr[29:7] == 2'd2);
	slave_sel[3] = (shared_adr[29:22] == 5'd16);
	slave_sel[4] = (shared_adr[29:26] == 2'd3);
	slave_sel[5] = (shared_adr[29:20] == 8'd152);
	slave_sel[6] = (shared_adr[29:14] == 16'd61440);
end
assign mgmtsoc_vexriscv_debug_bus_adr = shared_adr;
assign mgmtsoc_vexriscv_debug_bus_dat_w = shared_dat_w;
assign mgmtsoc_vexriscv_debug_bus_sel = shared_sel;
assign mgmtsoc_vexriscv_debug_bus_stb = shared_stb;
assign mgmtsoc_vexriscv_debug_bus_we = shared_we;
assign mgmtsoc_vexriscv_debug_bus_cti = shared_cti;
assign mgmtsoc_vexriscv_debug_bus_bte = shared_bte;
assign dff_bus_adr = shared_adr;
assign dff_bus_dat_w = shared_dat_w;
assign dff_bus_sel = shared_sel;
assign dff_bus_stb = shared_stb;
assign dff_bus_we = shared_we;
assign dff_bus_cti = shared_cti;
assign dff_bus_bte = shared_bte;
assign dff2_bus_adr = shared_adr;
assign dff2_bus_dat_w = shared_dat_w;
assign dff2_bus_sel = shared_sel;
assign dff2_bus_stb = shared_stb;
assign dff2_bus_we = shared_we;
assign dff2_bus_cti = shared_cti;
assign dff2_bus_bte = shared_bte;
assign mgmtsoc_litespimmap_bus_adr = shared_adr;
assign mgmtsoc_litespimmap_bus_dat_w = shared_dat_w;
assign mgmtsoc_litespimmap_bus_sel = shared_sel;
assign mgmtsoc_litespimmap_bus_stb = shared_stb;
assign mgmtsoc_litespimmap_bus_we = shared_we;
assign mgmtsoc_litespimmap_bus_cti = shared_cti;
assign mgmtsoc_litespimmap_bus_bte = shared_bte;
assign mprj_adr = shared_adr;
assign mprj_dat_w = shared_dat_w;
assign mprj_sel = shared_sel;
assign mprj_stb = shared_stb;
assign mprj_we = shared_we;
assign mprj_cti = shared_cti;
assign mprj_bte = shared_bte;
assign hk_adr = shared_adr;
assign hk_dat_w = shared_dat_w;
assign hk_sel = shared_sel;
assign hk_stb = shared_stb;
assign hk_we = shared_we;
assign hk_cti = shared_cti;
assign hk_bte = shared_bte;
assign mgmtsoc_wishbone_adr = shared_adr;
assign mgmtsoc_wishbone_dat_w = shared_dat_w;
assign mgmtsoc_wishbone_sel = shared_sel;
assign mgmtsoc_wishbone_stb = shared_stb;
assign mgmtsoc_wishbone_we = shared_we;
assign mgmtsoc_wishbone_cti = shared_cti;
assign mgmtsoc_wishbone_bte = shared_bte;
assign mgmtsoc_vexriscv_debug_bus_cyc = (shared_cyc & slave_sel[0]);
assign dff_bus_cyc = (shared_cyc & slave_sel[1]);
assign dff2_bus_cyc = (shared_cyc & slave_sel[2]);
assign mgmtsoc_litespimmap_bus_cyc = (shared_cyc & slave_sel[3]);
assign mprj_cyc = (shared_cyc & slave_sel[4]);
assign hk_cyc = (shared_cyc & slave_sel[5]);
assign mgmtsoc_wishbone_cyc = (shared_cyc & slave_sel[6]);
always @(*) begin
	shared_ack = 1'd0;
	shared_ack = ((((((mgmtsoc_vexriscv_debug_bus_ack | dff_bus_ack) | dff2_bus_ack) | mgmtsoc_litespimmap_bus_ack) | mprj_ack) | hk_ack) | mgmtsoc_wishbone_ack);
	if (done) begin
		shared_ack = 1'd1;
	end
end
assign shared_err = ((((((mgmtsoc_vexriscv_debug_bus_err | dff_bus_err) | dff2_bus_err) | mgmtsoc_litespimmap_bus_err) | mprj_err) | hk_err) | mgmtsoc_wishbone_err);
always @(*) begin
	shared_dat_r = 32'd0;
	shared_dat_r = ((((((({32{slave_sel_r[0]}} & mgmtsoc_vexriscv_debug_bus_dat_r) | ({32{slave_sel_r[1]}} & dff_bus_dat_r)) | ({32{slave_sel_r[2]}} & dff2_bus_dat_r)) | ({32{slave_sel_r[3]}} & mgmtsoc_litespimmap_bus_dat_r)) | ({32{slave_sel_r[4]}} & mprj_dat_r)) | ({32{slave_sel_r[5]}} & hk_dat_r)) | ({32{slave_sel_r[6]}} & mgmtsoc_wishbone_dat_r));
	if (done) begin
		shared_dat_r = 32'd4294967295;
	end
end
assign wait_1 = ((shared_stb & shared_cyc) & (~shared_ack));
always @(*) begin
	error = 1'd0;
	if (done) begin
		error = 1'd1;
	end
end
assign done = (count == 1'd0);
assign csrbank0_sel = (interface0_bank_bus_adr[13:9] == 1'd0);
assign csrbank0_reset0_r = interface0_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank0_reset0_re = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank0_reset0_re = interface0_bank_bus_we;
	end
end
always @(*) begin
	csrbank0_reset0_we = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank0_reset0_we = (~interface0_bank_bus_we);
	end
end
assign csrbank0_scratch0_r = interface0_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank0_scratch0_we = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank0_scratch0_we = (~interface0_bank_bus_we);
	end
end
always @(*) begin
	csrbank0_scratch0_re = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank0_scratch0_re = interface0_bank_bus_we;
	end
end
assign csrbank0_bus_errors_r = interface0_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank0_bus_errors_re = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank0_bus_errors_re = interface0_bank_bus_we;
	end
end
always @(*) begin
	csrbank0_bus_errors_we = 1'd0;
	if ((csrbank0_sel & (interface0_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank0_bus_errors_we = (~interface0_bank_bus_we);
	end
end
always @(*) begin
	mgmtsoc_soc_rst = 1'd0;
	if (mgmtsoc_reset_re) begin
		mgmtsoc_soc_rst = mgmtsoc_reset_storage[0];
	end
end
assign mgmtsoc_cpu_rst = mgmtsoc_reset_storage[1];
assign csrbank0_reset0_w = mgmtsoc_reset_storage[1:0];
assign csrbank0_scratch0_w = mgmtsoc_scratch_storage[31:0];
assign csrbank0_bus_errors_w = mgmtsoc_bus_errors_status[31:0];
assign mgmtsoc_bus_errors_we = csrbank0_bus_errors_we;
assign csrbank1_sel = (interface1_bank_bus_adr[13:9] == 1'd1);
assign csrbank1_out0_r = interface1_bank_bus_dat_w[0];
always @(*) begin
	csrbank1_out0_we = 1'd0;
	if ((csrbank1_sel & (interface1_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank1_out0_we = (~interface1_bank_bus_we);
	end
end
always @(*) begin
	csrbank1_out0_re = 1'd0;
	if ((csrbank1_sel & (interface1_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank1_out0_re = interface1_bank_bus_we;
	end
end
assign csrbank1_out0_w = debug_mode_storage;
assign csrbank2_sel = (interface2_bank_bus_adr[13:9] == 2'd2);
assign csrbank2_out0_r = interface2_bank_bus_dat_w[0];
always @(*) begin
	csrbank2_out0_we = 1'd0;
	if ((csrbank2_sel & (interface2_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank2_out0_we = (~interface2_bank_bus_we);
	end
end
always @(*) begin
	csrbank2_out0_re = 1'd0;
	if ((csrbank2_sel & (interface2_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank2_out0_re = interface2_bank_bus_we;
	end
end
assign csrbank2_out0_w = debug_oeb_storage;
assign csrbank3_sel = (interface3_bank_bus_adr[13:9] == 2'd3);
assign csrbank3_mmap_dummy_bits0_r = interface3_bank_bus_dat_w[7:0];
always @(*) begin
	csrbank3_mmap_dummy_bits0_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank3_mmap_dummy_bits0_re = interface3_bank_bus_we;
	end
end
always @(*) begin
	csrbank3_mmap_dummy_bits0_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank3_mmap_dummy_bits0_we = (~interface3_bank_bus_we);
	end
end
assign csrbank3_master_cs0_r = interface3_bank_bus_dat_w[0];
always @(*) begin
	csrbank3_master_cs0_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank3_master_cs0_re = interface3_bank_bus_we;
	end
end
always @(*) begin
	csrbank3_master_cs0_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank3_master_cs0_we = (~interface3_bank_bus_we);
	end
end
assign csrbank3_master_phyconfig0_r = interface3_bank_bus_dat_w[23:0];
always @(*) begin
	csrbank3_master_phyconfig0_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank3_master_phyconfig0_we = (~interface3_bank_bus_we);
	end
end
always @(*) begin
	csrbank3_master_phyconfig0_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank3_master_phyconfig0_re = interface3_bank_bus_we;
	end
end
assign mgmtsoc_master_rxtx_r = interface3_bank_bus_dat_w[31:0];
always @(*) begin
	mgmtsoc_master_rxtx_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 2'd3))) begin
		mgmtsoc_master_rxtx_re = interface3_bank_bus_we;
	end
end
always @(*) begin
	mgmtsoc_master_rxtx_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 2'd3))) begin
		mgmtsoc_master_rxtx_we = (~interface3_bank_bus_we);
	end
end
assign csrbank3_master_status_r = interface3_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank3_master_status_re = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank3_master_status_re = interface3_bank_bus_we;
	end
end
always @(*) begin
	csrbank3_master_status_we = 1'd0;
	if ((csrbank3_sel & (interface3_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank3_master_status_we = (~interface3_bank_bus_we);
	end
end
assign csrbank3_mmap_dummy_bits0_w = mgmtsoc_litespimmap_storage[7:0];
assign csrbank3_master_cs0_w = mgmtsoc_master_cs_storage;
assign mgmtsoc_master_len = mgmtsoc_master_phyconfig_storage[7:0];
assign mgmtsoc_master_width = mgmtsoc_master_phyconfig_storage[11:8];
assign mgmtsoc_master_mask = mgmtsoc_master_phyconfig_storage[23:16];
assign csrbank3_master_phyconfig0_w = mgmtsoc_master_phyconfig_storage[23:0];
always @(*) begin
	mgmtsoc_master_status_status = 2'd0;
	mgmtsoc_master_status_status[0] = mgmtsoc_master_tx_ready;
	mgmtsoc_master_status_status[1] = mgmtsoc_master_rx_ready;
end
assign csrbank3_master_status_w = mgmtsoc_master_status_status[1:0];
assign mgmtsoc_master_status_we = csrbank3_master_status_we;
assign csrbank4_sel = (interface4_bank_bus_adr[13:9] == 3'd4);
assign csrbank4_clk_divisor0_r = interface4_bank_bus_dat_w[7:0];
always @(*) begin
	csrbank4_clk_divisor0_we = 1'd0;
	if ((csrbank4_sel & (interface4_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank4_clk_divisor0_we = (~interface4_bank_bus_we);
	end
end
always @(*) begin
	csrbank4_clk_divisor0_re = 1'd0;
	if ((csrbank4_sel & (interface4_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank4_clk_divisor0_re = interface4_bank_bus_we;
	end
end
assign csrbank4_clk_divisor0_w = mgmtsoc_litespisdrphycore_storage[7:0];
assign csrbank5_sel = (interface5_bank_bus_adr[13:9] == 3'd5);
assign csrbank5_mode10_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_mode10_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank5_mode10_we = (~interface5_bank_bus_we);
	end
end
always @(*) begin
	csrbank5_mode10_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank5_mode10_re = interface5_bank_bus_we;
	end
end
assign csrbank5_mode00_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_mode00_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank5_mode00_re = interface5_bank_bus_we;
	end
end
always @(*) begin
	csrbank5_mode00_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank5_mode00_we = (~interface5_bank_bus_we);
	end
end
assign csrbank5_ien0_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_ien0_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank5_ien0_we = (~interface5_bank_bus_we);
	end
end
always @(*) begin
	csrbank5_ien0_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank5_ien0_re = interface5_bank_bus_we;
	end
end
assign csrbank5_oe0_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_oe0_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank5_oe0_we = (~interface5_bank_bus_we);
	end
end
always @(*) begin
	csrbank5_oe0_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank5_oe0_re = interface5_bank_bus_we;
	end
end
assign csrbank5_in_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_in_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank5_in_re = interface5_bank_bus_we;
	end
end
always @(*) begin
	csrbank5_in_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank5_in_we = (~interface5_bank_bus_we);
	end
end
assign csrbank5_out0_r = interface5_bank_bus_dat_w[0];
always @(*) begin
	csrbank5_out0_we = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank5_out0_we = (~interface5_bank_bus_we);
	end
end
always @(*) begin
	csrbank5_out0_re = 1'd0;
	if ((csrbank5_sel & (interface5_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank5_out0_re = interface5_bank_bus_we;
	end
end
assign csrbank5_mode10_w = gpio_mode1_storage;
assign csrbank5_mode00_w = gpio_mode0_storage;
assign csrbank5_ien0_w = gpio_ien_storage;
assign csrbank5_oe0_w = gpio_oe_storage;
assign csrbank5_in_w = gpio_in_status;
assign gpio_in_we = csrbank5_in_we;
assign csrbank5_out0_w = gpio_out_storage;
assign csrbank6_sel = (interface6_bank_bus_adr[13:9] == 3'd6);
assign csrbank6_ien3_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_ien3_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank6_ien3_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_ien3_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank6_ien3_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_ien2_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_ien2_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank6_ien2_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_ien2_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank6_ien2_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_ien1_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_ien1_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank6_ien1_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_ien1_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank6_ien1_re = interface6_bank_bus_we;
	end
end
assign csrbank6_ien0_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_ien0_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank6_ien0_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_ien0_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank6_ien0_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_oe3_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_oe3_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank6_oe3_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_oe3_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank6_oe3_re = interface6_bank_bus_we;
	end
end
assign csrbank6_oe2_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_oe2_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank6_oe2_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_oe2_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank6_oe2_re = interface6_bank_bus_we;
	end
end
assign csrbank6_oe1_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_oe1_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank6_oe1_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_oe1_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank6_oe1_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_oe0_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_oe0_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank6_oe0_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_oe0_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank6_oe0_re = interface6_bank_bus_we;
	end
end
assign csrbank6_in3_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_in3_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd8))) begin
		csrbank6_in3_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_in3_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd8))) begin
		csrbank6_in3_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_in2_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_in2_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd9))) begin
		csrbank6_in2_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_in2_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd9))) begin
		csrbank6_in2_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_in1_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_in1_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd10))) begin
		csrbank6_in1_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_in1_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd10))) begin
		csrbank6_in1_re = interface6_bank_bus_we;
	end
end
assign csrbank6_in0_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_in0_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd11))) begin
		csrbank6_in0_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_in0_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd11))) begin
		csrbank6_in0_re = interface6_bank_bus_we;
	end
end
assign csrbank6_out3_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_out3_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd12))) begin
		csrbank6_out3_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_out3_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd12))) begin
		csrbank6_out3_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_out2_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_out2_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd13))) begin
		csrbank6_out2_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_out2_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd13))) begin
		csrbank6_out2_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_out1_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_out1_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd14))) begin
		csrbank6_out1_we = (~interface6_bank_bus_we);
	end
end
always @(*) begin
	csrbank6_out1_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd14))) begin
		csrbank6_out1_re = interface6_bank_bus_we;
	end
end
assign csrbank6_out0_r = interface6_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank6_out0_re = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd15))) begin
		csrbank6_out0_re = interface6_bank_bus_we;
	end
end
always @(*) begin
	csrbank6_out0_we = 1'd0;
	if ((csrbank6_sel & (interface6_bank_bus_adr[8:0] == 4'd15))) begin
		csrbank6_out0_we = (~interface6_bank_bus_we);
	end
end
assign csrbank6_ien3_w = la_ien_storage[127:96];
assign csrbank6_ien2_w = la_ien_storage[95:64];
assign csrbank6_ien1_w = la_ien_storage[63:32];
assign csrbank6_ien0_w = la_ien_storage[31:0];
assign csrbank6_oe3_w = la_oe_storage[127:96];
assign csrbank6_oe2_w = la_oe_storage[95:64];
assign csrbank6_oe1_w = la_oe_storage[63:32];
assign csrbank6_oe0_w = la_oe_storage[31:0];
assign csrbank6_in3_w = la_in_status[127:96];
assign csrbank6_in2_w = la_in_status[95:64];
assign csrbank6_in1_w = la_in_status[63:32];
assign csrbank6_in0_w = la_in_status[31:0];
assign la_in_we = csrbank6_in0_we;
assign csrbank6_out3_w = la_out_storage[127:96];
assign csrbank6_out2_w = la_out_storage[95:64];
assign csrbank6_out1_w = la_out_storage[63:32];
assign csrbank6_out0_w = la_out_storage[31:0];
assign csrbank7_sel = (interface7_bank_bus_adr[13:9] == 3'd7);
assign csrbank7_out0_r = interface7_bank_bus_dat_w[0];
always @(*) begin
	csrbank7_out0_re = 1'd0;
	if ((csrbank7_sel & (interface7_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank7_out0_re = interface7_bank_bus_we;
	end
end
always @(*) begin
	csrbank7_out0_we = 1'd0;
	if ((csrbank7_sel & (interface7_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank7_out0_we = (~interface7_bank_bus_we);
	end
end
assign csrbank7_out0_w = mprj_wb_iena_storage;
assign csrbank8_sel = (interface8_bank_bus_adr[13:9] == 4'd8);
assign csrbank8_out0_r = interface8_bank_bus_dat_w[0];
always @(*) begin
	csrbank8_out0_we = 1'd0;
	if ((csrbank8_sel & (interface8_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank8_out0_we = (~interface8_bank_bus_we);
	end
end
always @(*) begin
	csrbank8_out0_re = 1'd0;
	if ((csrbank8_sel & (interface8_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank8_out0_re = interface8_bank_bus_we;
	end
end
assign csrbank8_out0_w = spi_enabled_storage;
assign csrbank9_sel = (interface9_bank_bus_adr[13:9] == 4'd9);
assign csrbank9_control0_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
	csrbank9_control0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank9_control0_we = (~interface9_bank_bus_we);
	end
end
always @(*) begin
	csrbank9_control0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank9_control0_re = interface9_bank_bus_we;
	end
end
assign csrbank9_status_r = interface9_bank_bus_dat_w[0];
always @(*) begin
	csrbank9_status_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank9_status_re = interface9_bank_bus_we;
	end
end
always @(*) begin
	csrbank9_status_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank9_status_we = (~interface9_bank_bus_we);
	end
end
assign csrbank9_mosi0_r = interface9_bank_bus_dat_w[7:0];
always @(*) begin
	csrbank9_mosi0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank9_mosi0_re = interface9_bank_bus_we;
	end
end
always @(*) begin
	csrbank9_mosi0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank9_mosi0_we = (~interface9_bank_bus_we);
	end
end
assign csrbank9_miso_r = interface9_bank_bus_dat_w[7:0];
always @(*) begin
	csrbank9_miso_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank9_miso_we = (~interface9_bank_bus_we);
	end
end
always @(*) begin
	csrbank9_miso_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank9_miso_re = interface9_bank_bus_we;
	end
end
assign csrbank9_cs0_r = interface9_bank_bus_dat_w[16:0];
always @(*) begin
	csrbank9_cs0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank9_cs0_we = (~interface9_bank_bus_we);
	end
end
always @(*) begin
	csrbank9_cs0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank9_cs0_re = interface9_bank_bus_we;
	end
end
assign csrbank9_loopback0_r = interface9_bank_bus_dat_w[0];
always @(*) begin
	csrbank9_loopback0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank9_loopback0_re = interface9_bank_bus_we;
	end
end
always @(*) begin
	csrbank9_loopback0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank9_loopback0_we = (~interface9_bank_bus_we);
	end
end
assign csrbank9_clk_divider0_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
	csrbank9_clk_divider0_we = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank9_clk_divider0_we = (~interface9_bank_bus_we);
	end
end
always @(*) begin
	csrbank9_clk_divider0_re = 1'd0;
	if ((csrbank9_sel & (interface9_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank9_clk_divider0_re = interface9_bank_bus_we;
	end
end
always @(*) begin
	spi_master_start1 = 1'd0;
	if (spi_master_control_re) begin
		spi_master_start1 = spi_master_control_storage[0];
	end
end
assign spi_master_length1 = spi_master_control_storage[15:8];
assign csrbank9_control0_w = spi_master_control_storage[15:0];
assign spi_master_status_status = spi_master_done1;
assign csrbank9_status_w = spi_master_status_status;
assign spi_master_status_we = csrbank9_status_we;
assign csrbank9_mosi0_w = spi_master_mosi_storage[7:0];
assign csrbank9_miso_w = spi_master_miso_status[7:0];
assign spi_master_miso_we = csrbank9_miso_we;
assign spi_master_sel = spi_master_cs_storage[0];
assign spi_master_mode0 = spi_master_cs_storage[16];
assign csrbank9_cs0_w = spi_master_cs_storage[16:0];
assign spi_master_mode1 = spi_master_loopback_storage;
assign csrbank9_loopback0_w = spi_master_loopback_storage;
assign csrbank9_clk_divider0_w = spimaster_storage[15:0];
assign csrbank10_sel = (interface10_bank_bus_adr[13:9] == 4'd10);
assign csrbank10_load0_r = interface10_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank10_load0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank10_load0_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_load0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank10_load0_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_reload0_r = interface10_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank10_reload0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank10_reload0_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_reload0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank10_reload0_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_en0_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_en0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank10_en0_we = (~interface10_bank_bus_we);
	end
end
always @(*) begin
	csrbank10_en0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank10_en0_re = interface10_bank_bus_we;
	end
end
assign csrbank10_update_value0_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_update_value0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank10_update_value0_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_update_value0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank10_update_value0_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_value_r = interface10_bank_bus_dat_w[31:0];
always @(*) begin
	csrbank10_value_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank10_value_we = (~interface10_bank_bus_we);
	end
end
always @(*) begin
	csrbank10_value_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank10_value_re = interface10_bank_bus_we;
	end
end
assign csrbank10_ev_status_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_ev_status_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank10_ev_status_we = (~interface10_bank_bus_we);
	end
end
always @(*) begin
	csrbank10_ev_status_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank10_ev_status_re = interface10_bank_bus_we;
	end
end
assign csrbank10_ev_pending_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_ev_pending_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank10_ev_pending_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_ev_pending_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank10_ev_pending_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_ev_enable0_r = interface10_bank_bus_dat_w[0];
always @(*) begin
	csrbank10_ev_enable0_re = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank10_ev_enable0_re = interface10_bank_bus_we;
	end
end
always @(*) begin
	csrbank10_ev_enable0_we = 1'd0;
	if ((csrbank10_sel & (interface10_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank10_ev_enable0_we = (~interface10_bank_bus_we);
	end
end
assign csrbank10_load0_w = mgmtsoc_load_storage[31:0];
assign csrbank10_reload0_w = mgmtsoc_reload_storage[31:0];
assign csrbank10_en0_w = mgmtsoc_en_storage;
assign csrbank10_update_value0_w = mgmtsoc_update_value_storage;
assign csrbank10_value_w = mgmtsoc_value_status[31:0];
assign mgmtsoc_value_we = csrbank10_value_we;
assign mgmtsoc_status_status = mgmtsoc_zero0;
assign csrbank10_ev_status_w = mgmtsoc_status_status;
assign mgmtsoc_status_we = csrbank10_ev_status_we;
assign mgmtsoc_pending_status = mgmtsoc_zero1;
assign csrbank10_ev_pending_w = mgmtsoc_pending_status;
assign mgmtsoc_pending_we = csrbank10_ev_pending_we;
assign mgmtsoc_zero2 = mgmtsoc_enable_storage;
assign csrbank10_ev_enable0_w = mgmtsoc_enable_storage;
assign csrbank11_sel = (interface11_bank_bus_adr[13:9] == 4'd11);
assign uart_rxtx_r = interface11_bank_bus_dat_w[7:0];
always @(*) begin
	uart_rxtx_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 1'd0))) begin
		uart_rxtx_we = (~interface11_bank_bus_we);
	end
end
always @(*) begin
	uart_rxtx_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 1'd0))) begin
		uart_rxtx_re = interface11_bank_bus_we;
	end
end
assign csrbank11_txfull_r = interface11_bank_bus_dat_w[0];
always @(*) begin
	csrbank11_txfull_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank11_txfull_we = (~interface11_bank_bus_we);
	end
end
always @(*) begin
	csrbank11_txfull_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank11_txfull_re = interface11_bank_bus_we;
	end
end
assign csrbank11_rxempty_r = interface11_bank_bus_dat_w[0];
always @(*) begin
	csrbank11_rxempty_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank11_rxempty_we = (~interface11_bank_bus_we);
	end
end
always @(*) begin
	csrbank11_rxempty_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank11_rxempty_re = interface11_bank_bus_we;
	end
end
assign csrbank11_ev_status_r = interface11_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank11_ev_status_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank11_ev_status_re = interface11_bank_bus_we;
	end
end
always @(*) begin
	csrbank11_ev_status_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank11_ev_status_we = (~interface11_bank_bus_we);
	end
end
assign csrbank11_ev_pending_r = interface11_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank11_ev_pending_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank11_ev_pending_re = interface11_bank_bus_we;
	end
end
always @(*) begin
	csrbank11_ev_pending_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank11_ev_pending_we = (~interface11_bank_bus_we);
	end
end
assign csrbank11_ev_enable0_r = interface11_bank_bus_dat_w[1:0];
always @(*) begin
	csrbank11_ev_enable0_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank11_ev_enable0_we = (~interface11_bank_bus_we);
	end
end
always @(*) begin
	csrbank11_ev_enable0_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank11_ev_enable0_re = interface11_bank_bus_we;
	end
end
assign csrbank11_txempty_r = interface11_bank_bus_dat_w[0];
always @(*) begin
	csrbank11_txempty_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank11_txempty_re = interface11_bank_bus_we;
	end
end
always @(*) begin
	csrbank11_txempty_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd6))) begin
		csrbank11_txempty_we = (~interface11_bank_bus_we);
	end
end
assign csrbank11_rxfull_r = interface11_bank_bus_dat_w[0];
always @(*) begin
	csrbank11_rxfull_re = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank11_rxfull_re = interface11_bank_bus_we;
	end
end
always @(*) begin
	csrbank11_rxfull_we = 1'd0;
	if ((csrbank11_sel & (interface11_bank_bus_adr[8:0] == 3'd7))) begin
		csrbank11_rxfull_we = (~interface11_bank_bus_we);
	end
end
assign csrbank11_txfull_w = uart_txfull_status;
assign uart_txfull_we = csrbank11_txfull_we;
assign csrbank11_rxempty_w = uart_rxempty_status;
assign uart_rxempty_we = csrbank11_rxempty_we;
always @(*) begin
	uart_status_status = 2'd0;
	uart_status_status[0] = uart_tx0;
	uart_status_status[1] = uart_rx0;
end
assign csrbank11_ev_status_w = uart_status_status[1:0];
assign uart_status_we = csrbank11_ev_status_we;
always @(*) begin
	uart_pending_status = 2'd0;
	uart_pending_status[0] = uart_tx1;
	uart_pending_status[1] = uart_rx1;
end
assign csrbank11_ev_pending_w = uart_pending_status[1:0];
assign uart_pending_we = csrbank11_ev_pending_we;
assign uart_tx2 = uart_enable_storage[0];
assign uart_rx2 = uart_enable_storage[1];
assign csrbank11_ev_enable0_w = uart_enable_storage[1:0];
assign csrbank11_txempty_w = uart_txempty_status;
assign uart_txempty_we = csrbank11_txempty_we;
assign csrbank11_rxfull_w = uart_rxfull_status;
assign uart_rxfull_we = csrbank11_rxfull_we;
assign csrbank12_sel = (interface12_bank_bus_adr[13:9] == 4'd12);
assign csrbank12_out0_r = interface12_bank_bus_dat_w[0];
always @(*) begin
	csrbank12_out0_we = 1'd0;
	if ((csrbank12_sel & (interface12_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank12_out0_we = (~interface12_bank_bus_we);
	end
end
always @(*) begin
	csrbank12_out0_re = 1'd0;
	if ((csrbank12_sel & (interface12_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank12_out0_re = interface12_bank_bus_we;
	end
end
assign csrbank12_out0_w = uart_enabled_storage;
assign csrbank13_sel = (interface13_bank_bus_adr[13:9] == 4'd13);
assign csrbank13_in_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_in_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank13_in_we = (~interface13_bank_bus_we);
	end
end
always @(*) begin
	csrbank13_in_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank13_in_re = interface13_bank_bus_we;
	end
end
assign csrbank13_mode0_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_mode0_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank13_mode0_we = (~interface13_bank_bus_we);
	end
end
always @(*) begin
	csrbank13_mode0_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank13_mode0_re = interface13_bank_bus_we;
	end
end
assign csrbank13_edge0_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_edge0_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank13_edge0_re = interface13_bank_bus_we;
	end
end
always @(*) begin
	csrbank13_edge0_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank13_edge0_we = (~interface13_bank_bus_we);
	end
end
assign csrbank13_ev_status_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_ev_status_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank13_ev_status_we = (~interface13_bank_bus_we);
	end
end
always @(*) begin
	csrbank13_ev_status_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank13_ev_status_re = interface13_bank_bus_we;
	end
end
assign csrbank13_ev_pending_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_ev_pending_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank13_ev_pending_we = (~interface13_bank_bus_we);
	end
end
always @(*) begin
	csrbank13_ev_pending_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank13_ev_pending_re = interface13_bank_bus_we;
	end
end
assign csrbank13_ev_enable0_r = interface13_bank_bus_dat_w[0];
always @(*) begin
	csrbank13_ev_enable0_re = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank13_ev_enable0_re = interface13_bank_bus_we;
	end
end
always @(*) begin
	csrbank13_ev_enable0_we = 1'd0;
	if ((csrbank13_sel & (interface13_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank13_ev_enable0_we = (~interface13_bank_bus_we);
	end
end
assign csrbank13_in_w = gpioin0_in_status;
assign gpioin0_in_we = csrbank13_in_we;
assign csrbank13_mode0_w = gpioin0_gpioin0_mode_storage;
assign csrbank13_edge0_w = gpioin0_gpioin0_edge_storage;
assign gpioin0_status_status = gpioin0_i00;
assign csrbank13_ev_status_w = gpioin0_status_status;
assign gpioin0_status_we = csrbank13_ev_status_we;
assign gpioin0_pending_status = gpioin0_i01;
assign csrbank13_ev_pending_w = gpioin0_pending_status;
assign gpioin0_pending_we = csrbank13_ev_pending_we;
assign gpioin0_i02 = gpioin0_enable_storage;
assign csrbank13_ev_enable0_w = gpioin0_enable_storage;
assign csrbank14_sel = (interface14_bank_bus_adr[13:9] == 4'd14);
assign csrbank14_in_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_in_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank14_in_we = (~interface14_bank_bus_we);
	end
end
always @(*) begin
	csrbank14_in_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank14_in_re = interface14_bank_bus_we;
	end
end
assign csrbank14_mode0_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_mode0_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank14_mode0_re = interface14_bank_bus_we;
	end
end
always @(*) begin
	csrbank14_mode0_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank14_mode0_we = (~interface14_bank_bus_we);
	end
end
assign csrbank14_edge0_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_edge0_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank14_edge0_re = interface14_bank_bus_we;
	end
end
always @(*) begin
	csrbank14_edge0_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank14_edge0_we = (~interface14_bank_bus_we);
	end
end
assign csrbank14_ev_status_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_ev_status_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank14_ev_status_we = (~interface14_bank_bus_we);
	end
end
always @(*) begin
	csrbank14_ev_status_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank14_ev_status_re = interface14_bank_bus_we;
	end
end
assign csrbank14_ev_pending_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_ev_pending_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank14_ev_pending_re = interface14_bank_bus_we;
	end
end
always @(*) begin
	csrbank14_ev_pending_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank14_ev_pending_we = (~interface14_bank_bus_we);
	end
end
assign csrbank14_ev_enable0_r = interface14_bank_bus_dat_w[0];
always @(*) begin
	csrbank14_ev_enable0_re = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank14_ev_enable0_re = interface14_bank_bus_we;
	end
end
always @(*) begin
	csrbank14_ev_enable0_we = 1'd0;
	if ((csrbank14_sel & (interface14_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank14_ev_enable0_we = (~interface14_bank_bus_we);
	end
end
assign csrbank14_in_w = gpioin1_in_status;
assign gpioin1_in_we = csrbank14_in_we;
assign csrbank14_mode0_w = gpioin1_gpioin1_mode_storage;
assign csrbank14_edge0_w = gpioin1_gpioin1_edge_storage;
assign gpioin1_status_status = gpioin1_i00;
assign csrbank14_ev_status_w = gpioin1_status_status;
assign gpioin1_status_we = csrbank14_ev_status_we;
assign gpioin1_pending_status = gpioin1_i01;
assign csrbank14_ev_pending_w = gpioin1_pending_status;
assign gpioin1_pending_we = csrbank14_ev_pending_we;
assign gpioin1_i02 = gpioin1_enable_storage;
assign csrbank14_ev_enable0_w = gpioin1_enable_storage;
assign csrbank15_sel = (interface15_bank_bus_adr[13:9] == 4'd15);
assign csrbank15_in_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_in_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank15_in_we = (~interface15_bank_bus_we);
	end
end
always @(*) begin
	csrbank15_in_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank15_in_re = interface15_bank_bus_we;
	end
end
assign csrbank15_mode0_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_mode0_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank15_mode0_re = interface15_bank_bus_we;
	end
end
always @(*) begin
	csrbank15_mode0_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank15_mode0_we = (~interface15_bank_bus_we);
	end
end
assign csrbank15_edge0_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_edge0_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank15_edge0_we = (~interface15_bank_bus_we);
	end
end
always @(*) begin
	csrbank15_edge0_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank15_edge0_re = interface15_bank_bus_we;
	end
end
assign csrbank15_ev_status_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_ev_status_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank15_ev_status_we = (~interface15_bank_bus_we);
	end
end
always @(*) begin
	csrbank15_ev_status_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank15_ev_status_re = interface15_bank_bus_we;
	end
end
assign csrbank15_ev_pending_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_ev_pending_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank15_ev_pending_re = interface15_bank_bus_we;
	end
end
always @(*) begin
	csrbank15_ev_pending_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank15_ev_pending_we = (~interface15_bank_bus_we);
	end
end
assign csrbank15_ev_enable0_r = interface15_bank_bus_dat_w[0];
always @(*) begin
	csrbank15_ev_enable0_we = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank15_ev_enable0_we = (~interface15_bank_bus_we);
	end
end
always @(*) begin
	csrbank15_ev_enable0_re = 1'd0;
	if ((csrbank15_sel & (interface15_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank15_ev_enable0_re = interface15_bank_bus_we;
	end
end
assign csrbank15_in_w = gpioin2_in_status;
assign gpioin2_in_we = csrbank15_in_we;
assign csrbank15_mode0_w = gpioin2_gpioin2_mode_storage;
assign csrbank15_edge0_w = gpioin2_gpioin2_edge_storage;
assign gpioin2_status_status = gpioin2_i00;
assign csrbank15_ev_status_w = gpioin2_status_status;
assign gpioin2_status_we = csrbank15_ev_status_we;
assign gpioin2_pending_status = gpioin2_i01;
assign csrbank15_ev_pending_w = gpioin2_pending_status;
assign gpioin2_pending_we = csrbank15_ev_pending_we;
assign gpioin2_i02 = gpioin2_enable_storage;
assign csrbank15_ev_enable0_w = gpioin2_enable_storage;
assign csrbank16_sel = (interface16_bank_bus_adr[13:9] == 5'd16);
assign csrbank16_in_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_in_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank16_in_re = interface16_bank_bus_we;
	end
end
always @(*) begin
	csrbank16_in_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank16_in_we = (~interface16_bank_bus_we);
	end
end
assign csrbank16_mode0_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_mode0_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank16_mode0_re = interface16_bank_bus_we;
	end
end
always @(*) begin
	csrbank16_mode0_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank16_mode0_we = (~interface16_bank_bus_we);
	end
end
assign csrbank16_edge0_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_edge0_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank16_edge0_we = (~interface16_bank_bus_we);
	end
end
always @(*) begin
	csrbank16_edge0_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank16_edge0_re = interface16_bank_bus_we;
	end
end
assign csrbank16_ev_status_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_ev_status_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank16_ev_status_re = interface16_bank_bus_we;
	end
end
always @(*) begin
	csrbank16_ev_status_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank16_ev_status_we = (~interface16_bank_bus_we);
	end
end
assign csrbank16_ev_pending_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_ev_pending_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank16_ev_pending_re = interface16_bank_bus_we;
	end
end
always @(*) begin
	csrbank16_ev_pending_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank16_ev_pending_we = (~interface16_bank_bus_we);
	end
end
assign csrbank16_ev_enable0_r = interface16_bank_bus_dat_w[0];
always @(*) begin
	csrbank16_ev_enable0_we = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank16_ev_enable0_we = (~interface16_bank_bus_we);
	end
end
always @(*) begin
	csrbank16_ev_enable0_re = 1'd0;
	if ((csrbank16_sel & (interface16_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank16_ev_enable0_re = interface16_bank_bus_we;
	end
end
assign csrbank16_in_w = gpioin3_in_status;
assign gpioin3_in_we = csrbank16_in_we;
assign csrbank16_mode0_w = gpioin3_gpioin3_mode_storage;
assign csrbank16_edge0_w = gpioin3_gpioin3_edge_storage;
assign gpioin3_status_status = gpioin3_i00;
assign csrbank16_ev_status_w = gpioin3_status_status;
assign gpioin3_status_we = csrbank16_ev_status_we;
assign gpioin3_pending_status = gpioin3_i01;
assign csrbank16_ev_pending_w = gpioin3_pending_status;
assign gpioin3_pending_we = csrbank16_ev_pending_we;
assign gpioin3_i02 = gpioin3_enable_storage;
assign csrbank16_ev_enable0_w = gpioin3_enable_storage;
assign csrbank17_sel = (interface17_bank_bus_adr[13:9] == 5'd17);
assign csrbank17_in_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_in_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank17_in_re = interface17_bank_bus_we;
	end
end
always @(*) begin
	csrbank17_in_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank17_in_we = (~interface17_bank_bus_we);
	end
end
assign csrbank17_mode0_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_mode0_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank17_mode0_re = interface17_bank_bus_we;
	end
end
always @(*) begin
	csrbank17_mode0_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank17_mode0_we = (~interface17_bank_bus_we);
	end
end
assign csrbank17_edge0_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_edge0_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank17_edge0_we = (~interface17_bank_bus_we);
	end
end
always @(*) begin
	csrbank17_edge0_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank17_edge0_re = interface17_bank_bus_we;
	end
end
assign csrbank17_ev_status_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_ev_status_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank17_ev_status_re = interface17_bank_bus_we;
	end
end
always @(*) begin
	csrbank17_ev_status_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank17_ev_status_we = (~interface17_bank_bus_we);
	end
end
assign csrbank17_ev_pending_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_ev_pending_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank17_ev_pending_re = interface17_bank_bus_we;
	end
end
always @(*) begin
	csrbank17_ev_pending_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank17_ev_pending_we = (~interface17_bank_bus_we);
	end
end
assign csrbank17_ev_enable0_r = interface17_bank_bus_dat_w[0];
always @(*) begin
	csrbank17_ev_enable0_we = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank17_ev_enable0_we = (~interface17_bank_bus_we);
	end
end
always @(*) begin
	csrbank17_ev_enable0_re = 1'd0;
	if ((csrbank17_sel & (interface17_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank17_ev_enable0_re = interface17_bank_bus_we;
	end
end
assign csrbank17_in_w = gpioin4_in_status;
assign gpioin4_in_we = csrbank17_in_we;
assign csrbank17_mode0_w = gpioin4_gpioin4_mode_storage;
assign csrbank17_edge0_w = gpioin4_gpioin4_edge_storage;
assign gpioin4_status_status = gpioin4_i00;
assign csrbank17_ev_status_w = gpioin4_status_status;
assign gpioin4_status_we = csrbank17_ev_status_we;
assign gpioin4_pending_status = gpioin4_i01;
assign csrbank17_ev_pending_w = gpioin4_pending_status;
assign gpioin4_pending_we = csrbank17_ev_pending_we;
assign gpioin4_i02 = gpioin4_enable_storage;
assign csrbank17_ev_enable0_w = gpioin4_enable_storage;
assign csrbank18_sel = (interface18_bank_bus_adr[13:9] == 5'd18);
assign csrbank18_in_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_in_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank18_in_re = interface18_bank_bus_we;
	end
end
always @(*) begin
	csrbank18_in_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank18_in_we = (~interface18_bank_bus_we);
	end
end
assign csrbank18_mode0_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_mode0_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank18_mode0_we = (~interface18_bank_bus_we);
	end
end
always @(*) begin
	csrbank18_mode0_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 1'd1))) begin
		csrbank18_mode0_re = interface18_bank_bus_we;
	end
end
assign csrbank18_edge0_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_edge0_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank18_edge0_we = (~interface18_bank_bus_we);
	end
end
always @(*) begin
	csrbank18_edge0_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 2'd2))) begin
		csrbank18_edge0_re = interface18_bank_bus_we;
	end
end
assign csrbank18_ev_status_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_ev_status_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank18_ev_status_re = interface18_bank_bus_we;
	end
end
always @(*) begin
	csrbank18_ev_status_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 2'd3))) begin
		csrbank18_ev_status_we = (~interface18_bank_bus_we);
	end
end
assign csrbank18_ev_pending_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_ev_pending_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank18_ev_pending_we = (~interface18_bank_bus_we);
	end
end
always @(*) begin
	csrbank18_ev_pending_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 3'd4))) begin
		csrbank18_ev_pending_re = interface18_bank_bus_we;
	end
end
assign csrbank18_ev_enable0_r = interface18_bank_bus_dat_w[0];
always @(*) begin
	csrbank18_ev_enable0_we = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank18_ev_enable0_we = (~interface18_bank_bus_we);
	end
end
always @(*) begin
	csrbank18_ev_enable0_re = 1'd0;
	if ((csrbank18_sel & (interface18_bank_bus_adr[8:0] == 3'd5))) begin
		csrbank18_ev_enable0_re = interface18_bank_bus_we;
	end
end
assign csrbank18_in_w = gpioin5_in_status;
assign gpioin5_in_we = csrbank18_in_we;
assign csrbank18_mode0_w = gpioin5_gpioin5_mode_storage;
assign csrbank18_edge0_w = gpioin5_gpioin5_edge_storage;
assign gpioin5_status_status = gpioin5_i00;
assign csrbank18_ev_status_w = gpioin5_status_status;
assign gpioin5_status_we = csrbank18_ev_status_we;
assign gpioin5_pending_status = gpioin5_i01;
assign csrbank18_ev_pending_w = gpioin5_pending_status;
assign gpioin5_pending_we = csrbank18_ev_pending_we;
assign gpioin5_i02 = gpioin5_enable_storage;
assign csrbank18_ev_enable0_w = gpioin5_enable_storage;
assign csrbank19_sel = (interface19_bank_bus_adr[13:9] == 5'd19);
assign csrbank19_out0_r = interface19_bank_bus_dat_w[2:0];
always @(*) begin
	csrbank19_out0_re = 1'd0;
	if ((csrbank19_sel & (interface19_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank19_out0_re = interface19_bank_bus_we;
	end
end
always @(*) begin
	csrbank19_out0_we = 1'd0;
	if ((csrbank19_sel & (interface19_bank_bus_adr[8:0] == 1'd0))) begin
		csrbank19_out0_we = (~interface19_bank_bus_we);
	end
end
assign csrbank19_out0_w = user_irq_ena_storage[2:0];
assign csr_interconnect_adr = mgmtsoc_adr;
assign csr_interconnect_we = mgmtsoc_we;
assign csr_interconnect_dat_w = mgmtsoc_dat_w;
assign mgmtsoc_dat_r = csr_interconnect_dat_r;
assign interface0_bank_bus_adr = csr_interconnect_adr;
assign interface1_bank_bus_adr = csr_interconnect_adr;
assign interface2_bank_bus_adr = csr_interconnect_adr;
assign interface3_bank_bus_adr = csr_interconnect_adr;
assign interface4_bank_bus_adr = csr_interconnect_adr;
assign interface5_bank_bus_adr = csr_interconnect_adr;
assign interface6_bank_bus_adr = csr_interconnect_adr;
assign interface7_bank_bus_adr = csr_interconnect_adr;
assign interface8_bank_bus_adr = csr_interconnect_adr;
assign interface9_bank_bus_adr = csr_interconnect_adr;
assign interface10_bank_bus_adr = csr_interconnect_adr;
assign interface11_bank_bus_adr = csr_interconnect_adr;
assign interface12_bank_bus_adr = csr_interconnect_adr;
assign interface13_bank_bus_adr = csr_interconnect_adr;
assign interface14_bank_bus_adr = csr_interconnect_adr;
assign interface15_bank_bus_adr = csr_interconnect_adr;
assign interface16_bank_bus_adr = csr_interconnect_adr;
assign interface17_bank_bus_adr = csr_interconnect_adr;
assign interface18_bank_bus_adr = csr_interconnect_adr;
assign interface19_bank_bus_adr = csr_interconnect_adr;
assign interface0_bank_bus_we = csr_interconnect_we;
assign interface1_bank_bus_we = csr_interconnect_we;
assign interface2_bank_bus_we = csr_interconnect_we;
assign interface3_bank_bus_we = csr_interconnect_we;
assign interface4_bank_bus_we = csr_interconnect_we;
assign interface5_bank_bus_we = csr_interconnect_we;
assign interface6_bank_bus_we = csr_interconnect_we;
assign interface7_bank_bus_we = csr_interconnect_we;
assign interface8_bank_bus_we = csr_interconnect_we;
assign interface9_bank_bus_we = csr_interconnect_we;
assign interface10_bank_bus_we = csr_interconnect_we;
assign interface11_bank_bus_we = csr_interconnect_we;
assign interface12_bank_bus_we = csr_interconnect_we;
assign interface13_bank_bus_we = csr_interconnect_we;
assign interface14_bank_bus_we = csr_interconnect_we;
assign interface15_bank_bus_we = csr_interconnect_we;
assign interface16_bank_bus_we = csr_interconnect_we;
assign interface17_bank_bus_we = csr_interconnect_we;
assign interface18_bank_bus_we = csr_interconnect_we;
assign interface19_bank_bus_we = csr_interconnect_we;
assign interface0_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface1_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface2_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface3_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface4_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface5_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface6_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface7_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface8_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface9_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface10_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface11_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface12_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface13_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface14_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface15_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface16_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface17_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface18_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface19_bank_bus_dat_w = csr_interconnect_dat_w;
assign csr_interconnect_dat_r = (((((((((((((((((((interface0_bank_bus_dat_r | interface1_bank_bus_dat_r) | interface2_bank_bus_dat_r) | interface3_bank_bus_dat_r) | interface4_bank_bus_dat_r) | interface5_bank_bus_dat_r) | interface6_bank_bus_dat_r) | interface7_bank_bus_dat_r) | interface8_bank_bus_dat_r) | interface9_bank_bus_dat_r) | interface10_bank_bus_dat_r) | interface11_bank_bus_dat_r) | interface12_bank_bus_dat_r) | interface13_bank_bus_dat_r) | interface14_bank_bus_dat_r) | interface15_bank_bus_dat_r) | interface16_bank_bus_dat_r) | interface17_bank_bus_dat_r) | interface18_bank_bus_dat_r) | interface19_bank_bus_dat_r);
always @(*) begin
	comb_array_muxed0 = 30'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed0 = mgmtsoc_ibus_ibus_adr;
		end
		1'd1: begin
			comb_array_muxed0 = mgmtsoc_dbus_dbus_adr;
		end
		default: begin
			comb_array_muxed0 = dbg_uart_wishbone_adr;
		end
	endcase
end
always @(*) begin
	comb_array_muxed1 = 32'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed1 = mgmtsoc_ibus_ibus_dat_w;
		end
		1'd1: begin
			comb_array_muxed1 = mgmtsoc_dbus_dbus_dat_w;
		end
		default: begin
			comb_array_muxed1 = dbg_uart_wishbone_dat_w;
		end
	endcase
end
always @(*) begin
	comb_array_muxed2 = 4'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed2 = mgmtsoc_ibus_ibus_sel;
		end
		1'd1: begin
			comb_array_muxed2 = mgmtsoc_dbus_dbus_sel;
		end
		default: begin
			comb_array_muxed2 = dbg_uart_wishbone_sel;
		end
	endcase
end
always @(*) begin
	comb_array_muxed3 = 1'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed3 = mgmtsoc_ibus_ibus_cyc;
		end
		1'd1: begin
			comb_array_muxed3 = mgmtsoc_dbus_dbus_cyc;
		end
		default: begin
			comb_array_muxed3 = dbg_uart_wishbone_cyc;
		end
	endcase
end
always @(*) begin
	comb_array_muxed4 = 1'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed4 = mgmtsoc_ibus_ibus_stb;
		end
		1'd1: begin
			comb_array_muxed4 = mgmtsoc_dbus_dbus_stb;
		end
		default: begin
			comb_array_muxed4 = dbg_uart_wishbone_stb;
		end
	endcase
end
always @(*) begin
	comb_array_muxed5 = 1'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed5 = mgmtsoc_ibus_ibus_we;
		end
		1'd1: begin
			comb_array_muxed5 = mgmtsoc_dbus_dbus_we;
		end
		default: begin
			comb_array_muxed5 = dbg_uart_wishbone_we;
		end
	endcase
end
always @(*) begin
	comb_array_muxed6 = 3'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed6 = mgmtsoc_ibus_ibus_cti;
		end
		1'd1: begin
			comb_array_muxed6 = mgmtsoc_dbus_dbus_cti;
		end
		default: begin
			comb_array_muxed6 = dbg_uart_wishbone_cti;
		end
	endcase
end
always @(*) begin
	comb_array_muxed7 = 2'd0;
	case (grant)
		1'd0: begin
			comb_array_muxed7 = mgmtsoc_ibus_ibus_bte;
		end
		1'd1: begin
			comb_array_muxed7 = mgmtsoc_dbus_dbus_bte;
		end
		default: begin
			comb_array_muxed7 = dbg_uart_wishbone_bte;
		end
	endcase
end
always @(*) begin
	sync_array_muxed = 1'd0;
	case (spi_master_mosi_sel)
		1'd0: begin
			sync_array_muxed = spi_master_mosi_data[0];
		end
		1'd1: begin
			sync_array_muxed = spi_master_mosi_data[1];
		end
		2'd2: begin
			sync_array_muxed = spi_master_mosi_data[2];
		end
		2'd3: begin
			sync_array_muxed = spi_master_mosi_data[3];
		end
		3'd4: begin
			sync_array_muxed = spi_master_mosi_data[4];
		end
		3'd5: begin
			sync_array_muxed = spi_master_mosi_data[5];
		end
		3'd6: begin
			sync_array_muxed = spi_master_mosi_data[6];
		end
		default: begin
			sync_array_muxed = spi_master_mosi_data[7];
		end
	endcase
end
assign sdrio_clk = sys_clk;
assign sdrio_clk_1 = sys_clk;
assign sdrio_clk_2 = sys_clk;
assign sdrio_clk_3 = sys_clk;
assign uart_phy_rx_rx = multiregimpl0_regs1;
assign dbg_uart_rx_rx = multiregimpl1_regs1;
assign gpio_in_status = multiregimpl2_regs1;
always @(*) begin
	la_in_status = 128'd0;
	la_in_status[0] = multiregimpl3_regs1;
	la_in_status[1] = multiregimpl4_regs1;
	la_in_status[2] = multiregimpl5_regs1;
	la_in_status[3] = multiregimpl6_regs1;
	la_in_status[4] = multiregimpl7_regs1;
	la_in_status[5] = multiregimpl8_regs1;
	la_in_status[6] = multiregimpl9_regs1;
	la_in_status[7] = multiregimpl10_regs1;
	la_in_status[8] = multiregimpl11_regs1;
	la_in_status[9] = multiregimpl12_regs1;
	la_in_status[10] = multiregimpl13_regs1;
	la_in_status[11] = multiregimpl14_regs1;
	la_in_status[12] = multiregimpl15_regs1;
	la_in_status[13] = multiregimpl16_regs1;
	la_in_status[14] = multiregimpl17_regs1;
	la_in_status[15] = multiregimpl18_regs1;
	la_in_status[16] = multiregimpl19_regs1;
	la_in_status[17] = multiregimpl20_regs1;
	la_in_status[18] = multiregimpl21_regs1;
	la_in_status[19] = multiregimpl22_regs1;
	la_in_status[20] = multiregimpl23_regs1;
	la_in_status[21] = multiregimpl24_regs1;
	la_in_status[22] = multiregimpl25_regs1;
	la_in_status[23] = multiregimpl26_regs1;
	la_in_status[24] = multiregimpl27_regs1;
	la_in_status[25] = multiregimpl28_regs1;
	la_in_status[26] = multiregimpl29_regs1;
	la_in_status[27] = multiregimpl30_regs1;
	la_in_status[28] = multiregimpl31_regs1;
	la_in_status[29] = multiregimpl32_regs1;
	la_in_status[30] = multiregimpl33_regs1;
	la_in_status[31] = multiregimpl34_regs1;
	la_in_status[32] = multiregimpl35_regs1;
	la_in_status[33] = multiregimpl36_regs1;
	la_in_status[34] = multiregimpl37_regs1;
	la_in_status[35] = multiregimpl38_regs1;
	la_in_status[36] = multiregimpl39_regs1;
	la_in_status[37] = multiregimpl40_regs1;
	la_in_status[38] = multiregimpl41_regs1;
	la_in_status[39] = multiregimpl42_regs1;
	la_in_status[40] = multiregimpl43_regs1;
	la_in_status[41] = multiregimpl44_regs1;
	la_in_status[42] = multiregimpl45_regs1;
	la_in_status[43] = multiregimpl46_regs1;
	la_in_status[44] = multiregimpl47_regs1;
	la_in_status[45] = multiregimpl48_regs1;
	la_in_status[46] = multiregimpl49_regs1;
	la_in_status[47] = multiregimpl50_regs1;
	la_in_status[48] = multiregimpl51_regs1;
	la_in_status[49] = multiregimpl52_regs1;
	la_in_status[50] = multiregimpl53_regs1;
	la_in_status[51] = multiregimpl54_regs1;
	la_in_status[52] = multiregimpl55_regs1;
	la_in_status[53] = multiregimpl56_regs1;
	la_in_status[54] = multiregimpl57_regs1;
	la_in_status[55] = multiregimpl58_regs1;
	la_in_status[56] = multiregimpl59_regs1;
	la_in_status[57] = multiregimpl60_regs1;
	la_in_status[58] = multiregimpl61_regs1;
	la_in_status[59] = multiregimpl62_regs1;
	la_in_status[60] = multiregimpl63_regs1;
	la_in_status[61] = multiregimpl64_regs1;
	la_in_status[62] = multiregimpl65_regs1;
	la_in_status[63] = multiregimpl66_regs1;
	la_in_status[64] = multiregimpl67_regs1;
	la_in_status[65] = multiregimpl68_regs1;
	la_in_status[66] = multiregimpl69_regs1;
	la_in_status[67] = multiregimpl70_regs1;
	la_in_status[68] = multiregimpl71_regs1;
	la_in_status[69] = multiregimpl72_regs1;
	la_in_status[70] = multiregimpl73_regs1;
	la_in_status[71] = multiregimpl74_regs1;
	la_in_status[72] = multiregimpl75_regs1;
	la_in_status[73] = multiregimpl76_regs1;
	la_in_status[74] = multiregimpl77_regs1;
	la_in_status[75] = multiregimpl78_regs1;
	la_in_status[76] = multiregimpl79_regs1;
	la_in_status[77] = multiregimpl80_regs1;
	la_in_status[78] = multiregimpl81_regs1;
	la_in_status[79] = multiregimpl82_regs1;
	la_in_status[80] = multiregimpl83_regs1;
	la_in_status[81] = multiregimpl84_regs1;
	la_in_status[82] = multiregimpl85_regs1;
	la_in_status[83] = multiregimpl86_regs1;
	la_in_status[84] = multiregimpl87_regs1;
	la_in_status[85] = multiregimpl88_regs1;
	la_in_status[86] = multiregimpl89_regs1;
	la_in_status[87] = multiregimpl90_regs1;
	la_in_status[88] = multiregimpl91_regs1;
	la_in_status[89] = multiregimpl92_regs1;
	la_in_status[90] = multiregimpl93_regs1;
	la_in_status[91] = multiregimpl94_regs1;
	la_in_status[92] = multiregimpl95_regs1;
	la_in_status[93] = multiregimpl96_regs1;
	la_in_status[94] = multiregimpl97_regs1;
	la_in_status[95] = multiregimpl98_regs1;
	la_in_status[96] = multiregimpl99_regs1;
	la_in_status[97] = multiregimpl100_regs1;
	la_in_status[98] = multiregimpl101_regs1;
	la_in_status[99] = multiregimpl102_regs1;
	la_in_status[100] = multiregimpl103_regs1;
	la_in_status[101] = multiregimpl104_regs1;
	la_in_status[102] = multiregimpl105_regs1;
	la_in_status[103] = multiregimpl106_regs1;
	la_in_status[104] = multiregimpl107_regs1;
	la_in_status[105] = multiregimpl108_regs1;
	la_in_status[106] = multiregimpl109_regs1;
	la_in_status[107] = multiregimpl110_regs1;
	la_in_status[108] = multiregimpl111_regs1;
	la_in_status[109] = multiregimpl112_regs1;
	la_in_status[110] = multiregimpl113_regs1;
	la_in_status[111] = multiregimpl114_regs1;
	la_in_status[112] = multiregimpl115_regs1;
	la_in_status[113] = multiregimpl116_regs1;
	la_in_status[114] = multiregimpl117_regs1;
	la_in_status[115] = multiregimpl118_regs1;
	la_in_status[116] = multiregimpl119_regs1;
	la_in_status[117] = multiregimpl120_regs1;
	la_in_status[118] = multiregimpl121_regs1;
	la_in_status[119] = multiregimpl122_regs1;
	la_in_status[120] = multiregimpl123_regs1;
	la_in_status[121] = multiregimpl124_regs1;
	la_in_status[122] = multiregimpl125_regs1;
	la_in_status[123] = multiregimpl126_regs1;
	la_in_status[124] = multiregimpl127_regs1;
	la_in_status[125] = multiregimpl128_regs1;
	la_in_status[126] = multiregimpl129_regs1;
	la_in_status[127] = multiregimpl130_regs1;
end
assign gpioin0_in_status = multiregimpl131_regs1;
assign gpioin1_in_status = multiregimpl132_regs1;
assign gpioin2_in_status = multiregimpl133_regs1;
assign gpioin3_in_status = multiregimpl134_regs1;
assign gpioin4_in_status = multiregimpl135_regs1;
assign gpioin5_in_status = multiregimpl136_regs1;

always @(posedge por_clk) begin
	int_rst <= core_rst;
end

always @(posedge sdrio_clk) begin
	flash_clk <= mgmtsoc_litespisdrphycore_clk;
	flash_io0_oeb <= (~mgmtsoc_litespisdrphycore_dq_oe);
	flash_io0_do <= mgmtsoc_litespisdrphycore_dq_o;
	mgmtsoc_litespisdrphycore_dq_i[1] <= flash_io1_di;
end

always @(posedge sys_clk) begin
	if ((mgmtsoc_bus_errors != 32'd4294967295)) begin
		if (mgmtsoc_bus_error) begin
			mgmtsoc_bus_errors <= (mgmtsoc_bus_errors + 1'd1);
		end
	end
	mgmtsoc_vexriscv_debug_bus_dat_r <= mgmtsoc_vexriscv_o_rsp_data;
	mgmtsoc_vexriscv_debug_reset <= (mgmtsoc_vexriscv_reset_debug_logic | sys_rst);
	if (((((mgmtsoc_vexriscv_debug_bus_stb & mgmtsoc_vexriscv_debug_bus_cyc) & (~mgmtsoc_vexriscv_transfer_in_progress)) & (~mgmtsoc_vexriscv_transfer_complete)) & (~mgmtsoc_vexriscv_transfer_wait_for_ack))) begin
		mgmtsoc_vexriscv_i_cmd_payload_data <= mgmtsoc_vexriscv_debug_bus_dat_w;
		mgmtsoc_vexriscv_i_cmd_payload_address <= ((mgmtsoc_vexriscv_debug_bus_adr[5:0] <<< 2'd2) | 1'd0);
		mgmtsoc_vexriscv_i_cmd_payload_wr <= mgmtsoc_vexriscv_debug_bus_we;
		mgmtsoc_vexriscv_i_cmd_valid <= 1'd1;
		mgmtsoc_vexriscv_transfer_in_progress <= 1'd1;
		mgmtsoc_vexriscv_transfer_complete <= 1'd0;
		mgmtsoc_vexriscv_debug_bus_ack <= 1'd0;
	end else begin
		if (mgmtsoc_vexriscv_transfer_in_progress) begin
			if (mgmtsoc_vexriscv_o_cmd_ready) begin
				mgmtsoc_vexriscv_i_cmd_valid <= 1'd0;
				mgmtsoc_vexriscv_i_cmd_payload_wr <= 1'd0;
				mgmtsoc_vexriscv_transfer_complete <= 1'd1;
				mgmtsoc_vexriscv_transfer_in_progress <= 1'd0;
			end
		end else begin
			if (mgmtsoc_vexriscv_transfer_complete) begin
				mgmtsoc_vexriscv_transfer_complete <= 1'd0;
				mgmtsoc_vexriscv_debug_bus_ack <= 1'd1;
				mgmtsoc_vexriscv_transfer_wait_for_ack <= 1'd1;
			end else begin
				if ((mgmtsoc_vexriscv_transfer_wait_for_ack & (~(mgmtsoc_vexriscv_debug_bus_stb & mgmtsoc_vexriscv_debug_bus_cyc)))) begin
					mgmtsoc_vexriscv_transfer_wait_for_ack <= 1'd0;
					mgmtsoc_vexriscv_debug_bus_ack <= 1'd0;
				end
			end
		end
	end
	if (mgmtsoc_vexriscv_o_resetOut) begin
		if ((mgmtsoc_ibus_ibus_cyc & mgmtsoc_ibus_ibus_stb)) begin
			mgmtsoc_vexriscv_ibus_err <= 1'd1;
		end else begin
			mgmtsoc_vexriscv_ibus_err <= 1'd0;
		end
		if ((mgmtsoc_dbus_dbus_cyc & mgmtsoc_dbus_dbus_stb)) begin
			mgmtsoc_vexriscv_dbus_err <= 1'd1;
		end else begin
			mgmtsoc_vexriscv_dbus_err <= 1'd0;
		end
		mgmtsoc_vexriscv_reset_debug_logic <= 1'd1;
	end else begin
		mgmtsoc_vexriscv_reset_debug_logic <= 1'd0;
	end
	if (mgmtsoc_en_storage) begin
		if ((mgmtsoc_value == 1'd0)) begin
			mgmtsoc_value <= mgmtsoc_reload_storage;
		end else begin
			mgmtsoc_value <= (mgmtsoc_value - 1'd1);
		end
	end else begin
		mgmtsoc_value <= mgmtsoc_load_storage;
	end
	if (mgmtsoc_update_value_re) begin
		mgmtsoc_value_status <= mgmtsoc_value;
	end
	if (mgmtsoc_zero_clear) begin
		mgmtsoc_zero_pending <= 1'd0;
	end
	mgmtsoc_zero_trigger_d <= mgmtsoc_zero_trigger;
	if ((mgmtsoc_zero_trigger & (~mgmtsoc_zero_trigger_d))) begin
		mgmtsoc_zero_pending <= 1'd1;
	end
	dff_bus_ack <= ((dff_bus_stb & dff_bus_cyc) & (~dff_bus_ack));
	dff2_bus_ack <= ((dff2_bus_stb & dff2_bus_cyc) & (~dff2_bus_ack));
	if (mgmtsoc_litespisdrphycore_sr_out_load) begin
		mgmtsoc_litespisdrphycore_sr_out <= (mgmtsoc_litespisdrphycore_sink_payload_data <<< (6'd32 - mgmtsoc_litespisdrphycore_sink_payload_len));
	end
	if (mgmtsoc_litespisdrphycore_sr_out_shift) begin
		case (mgmtsoc_litespisdrphycore_sink_payload_width)
			1'd1: begin
				mgmtsoc_litespisdrphycore_sr_out <= {mgmtsoc_litespisdrphycore_sr_out, mgmtsoc_litespisdrphycore0};
			end
			2'd2: begin
				mgmtsoc_litespisdrphycore_sr_out <= {mgmtsoc_litespisdrphycore_sr_out, mgmtsoc_litespisdrphycore1};
			end
			3'd4: begin
				mgmtsoc_litespisdrphycore_sr_out <= {mgmtsoc_litespisdrphycore_sr_out, mgmtsoc_litespisdrphycore2};
			end
			4'd8: begin
				mgmtsoc_litespisdrphycore_sr_out <= {mgmtsoc_litespisdrphycore_sr_out, mgmtsoc_litespisdrphycore3};
			end
		endcase
	end
	if (mgmtsoc_litespisdrphycore_sr_in_shift) begin
		case (mgmtsoc_litespisdrphycore_sink_payload_width)
			1'd1: begin
				mgmtsoc_litespisdrphycore_sr_in <= {mgmtsoc_litespisdrphycore_sr_in, mgmtsoc_litespisdrphycore_dq_i[1]};
			end
			2'd2: begin
				mgmtsoc_litespisdrphycore_sr_in <= {mgmtsoc_litespisdrphycore_sr_in, mgmtsoc_litespisdrphycore_dq_i[1:0]};
			end
			3'd4: begin
				mgmtsoc_litespisdrphycore_sr_in <= {mgmtsoc_litespisdrphycore_sr_in, mgmtsoc_litespisdrphycore_dq_i[1:0]};
			end
			4'd8: begin
				mgmtsoc_litespisdrphycore_sr_in <= {mgmtsoc_litespisdrphycore_sr_in, mgmtsoc_litespisdrphycore_dq_i[1:0]};
			end
		endcase
	end
	mgmtsoc_litespisdrphycore_posedge_reg <= mgmtsoc_litespisdrphycore_posedge;
	mgmtsoc_litespisdrphycore_posedge_reg2 <= mgmtsoc_litespisdrphycore_posedge_reg;
	if ((mgmtsoc_litespisdrphycore_en | mgmtsoc_litespisdrphycore_en_int)) begin
		if ((mgmtsoc_litespisdrphycore_cnt < mgmtsoc_litespisdrphycore_div)) begin
			mgmtsoc_litespisdrphycore_cnt <= (mgmtsoc_litespisdrphycore_cnt + 1'd1);
		end else begin
			mgmtsoc_litespisdrphycore_cnt <= 1'd0;
			mgmtsoc_litespisdrphycore_clk <= (~mgmtsoc_litespisdrphycore_clk);
		end
	end else begin
		mgmtsoc_litespisdrphycore_clk <= 1'd0;
		mgmtsoc_litespisdrphycore_cnt <= 1'd0;
	end
	if (mgmtsoc_litespisdrphycore_wait) begin
		if ((~mgmtsoc_litespisdrphycore_done)) begin
			mgmtsoc_litespisdrphycore_count <= (mgmtsoc_litespisdrphycore_count - 1'd1);
		end
	end else begin
		mgmtsoc_litespisdrphycore_count <= 4'd11;
	end
	litespiphy_state <= litespiphy_next_state;
	if (mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value_ce) begin
		mgmtsoc_litespisdrphycore_sr_cnt <= mgmtsoc_litespisdrphycore_sr_cnt_litespiphy_next_value;
	end
	case (litespi_grant)
		1'd0: begin
			if ((~litespi_request[0])) begin
				if (litespi_request[1]) begin
					litespi_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~litespi_request[1])) begin
				if (litespi_request[0]) begin
					litespi_grant <= 1'd0;
				end
			end
		end
	endcase
	if (mgmtsoc_litespimmap_wait) begin
		if ((~mgmtsoc_litespimmap_done)) begin
			mgmtsoc_litespimmap_count <= (mgmtsoc_litespimmap_count - 1'd1);
		end
	end else begin
		mgmtsoc_litespimmap_count <= 9'd256;
	end
	litespi_state <= litespi_next_state;
	if (mgmtsoc_litespimmap_burst_cs_litespi_next_value_ce0) begin
		mgmtsoc_litespimmap_burst_cs <= mgmtsoc_litespimmap_burst_cs_litespi_next_value0;
	end
	if (mgmtsoc_litespimmap_burst_adr_litespi_next_value_ce1) begin
		mgmtsoc_litespimmap_burst_adr <= mgmtsoc_litespimmap_burst_adr_litespi_next_value1;
	end
	if (((~mgmtsoc_master_tx_fifo_source_valid) | mgmtsoc_master_tx_fifo_source_ready)) begin
		mgmtsoc_master_tx_fifo_source_valid <= mgmtsoc_master_tx_fifo_sink_valid;
		mgmtsoc_master_tx_fifo_source_first <= mgmtsoc_master_tx_fifo_sink_first;
		mgmtsoc_master_tx_fifo_source_last <= mgmtsoc_master_tx_fifo_sink_last;
		mgmtsoc_master_tx_fifo_source_payload_data <= mgmtsoc_master_tx_fifo_sink_payload_data;
		mgmtsoc_master_tx_fifo_source_payload_len <= mgmtsoc_master_tx_fifo_sink_payload_len;
		mgmtsoc_master_tx_fifo_source_payload_width <= mgmtsoc_master_tx_fifo_sink_payload_width;
		mgmtsoc_master_tx_fifo_source_payload_mask <= mgmtsoc_master_tx_fifo_sink_payload_mask;
	end
	if (((~mgmtsoc_master_rx_fifo_source_valid) | mgmtsoc_master_rx_fifo_source_ready)) begin
		mgmtsoc_master_rx_fifo_source_valid <= mgmtsoc_master_rx_fifo_sink_valid;
		mgmtsoc_master_rx_fifo_source_first <= mgmtsoc_master_rx_fifo_sink_first;
		mgmtsoc_master_rx_fifo_source_last <= mgmtsoc_master_rx_fifo_sink_last;
		mgmtsoc_master_rx_fifo_source_payload_data <= mgmtsoc_master_rx_fifo_sink_payload_data;
	end
	spi_master_clk_divider1 <= (spi_master_clk_divider1 + 1'd1);
	if (spi_master_clk_rise) begin
		spi_clk <= spi_master_clk_enable;
	end else begin
		if (spi_master_clk_fall) begin
			spi_master_clk_divider1 <= 1'd0;
			spi_clk <= 1'd0;
		end
	end
	spi_cs_n <= (~(spi_master_cs & (spi_master_xfer_enable | (spi_master_cs_mode == 1'd1))));
	if (spi_master_mosi_latch) begin
		spi_master_mosi_data <= spi_master_mosi;
		spi_master_mosi_sel <= 3'd7;
	end else begin
		if (spi_master_clk_fall) begin
			if (spi_master_xfer_enable) begin
				spi_mosi <= sync_array_muxed;
			end
			spi_master_mosi_sel <= (spi_master_mosi_sel - 1'd1);
		end
	end
	if (spi_master_clk_rise) begin
		if (spi_master_loopback) begin
			spi_master_miso_data <= {spi_master_miso_data, spi_mosi};
		end else begin
			spi_master_miso_data <= {spi_master_miso_data, spi_miso};
		end
	end
	if (spi_master_miso_latch) begin
		spi_master_miso <= spi_master_miso_data;
	end
	spimaster_state <= spimaster_next_state;
	if (spi_master_count_spimaster_next_value_ce) begin
		spi_master_count <= spi_master_count_spimaster_next_value;
	end
	{uart_phy_tx_tick, uart_phy_tx_phase} <= 22'd4123168;
	if (uart_phy_tx_enable) begin
		{uart_phy_tx_tick, uart_phy_tx_phase} <= (uart_phy_tx_phase + 22'd4123168);
	end
	rs232phy_rs232phytx_state <= rs232phy_rs232phytx_next_state;
	if (uart_phy_tx_count_rs232phy_rs232phytx_next_value_ce0) begin
		uart_phy_tx_count <= uart_phy_tx_count_rs232phy_rs232phytx_next_value0;
	end
	if (sys_uart_tx_rs232phy_rs232phytx_next_value_ce1) begin
		sys_uart_tx <= sys_uart_tx_rs232phy_rs232phytx_next_value1;
	end
	if (uart_phy_tx_data_rs232phy_rs232phytx_next_value_ce2) begin
		uart_phy_tx_data <= uart_phy_tx_data_rs232phy_rs232phytx_next_value2;
	end
	uart_phy_rx_rx_d <= uart_phy_rx_rx;
	{uart_phy_rx_tick, uart_phy_rx_phase} <= 32'd2147483648;
	if (uart_phy_rx_enable) begin
		{uart_phy_rx_tick, uart_phy_rx_phase} <= (uart_phy_rx_phase + 22'd4123168);
	end
	rs232phy_rs232phyrx_state <= rs232phy_rs232phyrx_next_state;
	if (uart_phy_rx_count_rs232phy_rs232phyrx_next_value_ce0) begin
		uart_phy_rx_count <= uart_phy_rx_count_rs232phy_rs232phyrx_next_value0;
	end
	if (uart_phy_rx_data_rs232phy_rs232phyrx_next_value_ce1) begin
		uart_phy_rx_data <= uart_phy_rx_data_rs232phy_rs232phyrx_next_value1;
	end
	if (uart_tx_clear) begin
		uart_tx_pending <= 1'd0;
	end
	uart_tx_trigger_d <= uart_tx_trigger;
	if ((uart_tx_trigger & (~uart_tx_trigger_d))) begin
		uart_tx_pending <= 1'd1;
	end
	if (uart_rx_clear) begin
		uart_rx_pending <= 1'd0;
	end
	uart_rx_trigger_d <= uart_rx_trigger;
	if ((uart_rx_trigger & (~uart_rx_trigger_d))) begin
		uart_rx_pending <= 1'd1;
	end
	if (uart_tx_fifo_syncfifo_re) begin
		uart_tx_fifo_readable <= 1'd1;
	end else begin
		if (uart_tx_fifo_re) begin
			uart_tx_fifo_readable <= 1'd0;
		end
	end
	if (((uart_tx_fifo_syncfifo_we & uart_tx_fifo_syncfifo_writable) & (~uart_tx_fifo_replace))) begin
		uart_tx_fifo_produce <= (uart_tx_fifo_produce + 1'd1);
	end
	if (uart_tx_fifo_do_read) begin
		uart_tx_fifo_consume <= (uart_tx_fifo_consume + 1'd1);
	end
	if (((uart_tx_fifo_syncfifo_we & uart_tx_fifo_syncfifo_writable) & (~uart_tx_fifo_replace))) begin
		if ((~uart_tx_fifo_do_read)) begin
			uart_tx_fifo_level0 <= (uart_tx_fifo_level0 + 1'd1);
		end
	end else begin
		if (uart_tx_fifo_do_read) begin
			uart_tx_fifo_level0 <= (uart_tx_fifo_level0 - 1'd1);
		end
	end
	if (uart_rx_fifo_syncfifo_re) begin
		uart_rx_fifo_readable <= 1'd1;
	end else begin
		if (uart_rx_fifo_re) begin
			uart_rx_fifo_readable <= 1'd0;
		end
	end
	if (((uart_rx_fifo_syncfifo_we & uart_rx_fifo_syncfifo_writable) & (~uart_rx_fifo_replace))) begin
		uart_rx_fifo_produce <= (uart_rx_fifo_produce + 1'd1);
	end
	if (uart_rx_fifo_do_read) begin
		uart_rx_fifo_consume <= (uart_rx_fifo_consume + 1'd1);
	end
	if (((uart_rx_fifo_syncfifo_we & uart_rx_fifo_syncfifo_writable) & (~uart_rx_fifo_replace))) begin
		if ((~uart_rx_fifo_do_read)) begin
			uart_rx_fifo_level0 <= (uart_rx_fifo_level0 + 1'd1);
		end
	end else begin
		if (uart_rx_fifo_do_read) begin
			uart_rx_fifo_level0 <= (uart_rx_fifo_level0 - 1'd1);
		end
	end
	{dbg_uart_tx_tick, dbg_uart_tx_phase} <= 26'd49478023;
	if (dbg_uart_tx_enable) begin
		{dbg_uart_tx_tick, dbg_uart_tx_phase} <= (dbg_uart_tx_phase + 26'd49478023);
	end
	uartwishbonebridge_rs232phytx_state <= uartwishbonebridge_rs232phytx_next_state;
	if (dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value_ce0) begin
		dbg_uart_tx_count <= dbg_uart_tx_count_uartwishbonebridge_rs232phytx_next_value0;
	end
	if (dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value_ce1) begin
		dbg_uart_dbg_uart_tx <= dbg_uart_dbg_uart_tx_uartwishbonebridge_rs232phytx_next_value1;
	end
	if (dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value_ce2) begin
		dbg_uart_tx_data <= dbg_uart_tx_data_uartwishbonebridge_rs232phytx_next_value2;
	end
	dbg_uart_rx_rx_d <= dbg_uart_rx_rx;
	{dbg_uart_rx_tick, dbg_uart_rx_phase} <= 32'd2147483648;
	if (dbg_uart_rx_enable) begin
		{dbg_uart_rx_tick, dbg_uart_rx_phase} <= (dbg_uart_rx_phase + 26'd49478023);
	end
	uartwishbonebridge_rs232phyrx_state <= uartwishbonebridge_rs232phyrx_next_state;
	if (dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value_ce0) begin
		dbg_uart_rx_count <= dbg_uart_rx_count_uartwishbonebridge_rs232phyrx_next_value0;
	end
	if (dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value_ce1) begin
		dbg_uart_rx_data <= dbg_uart_rx_data_uartwishbonebridge_rs232phyrx_next_value1;
	end
	uartwishbonebridge_state <= uartwishbonebridge_next_state;
	if (dbg_uart_bytes_count_uartwishbonebridge_next_value_ce0) begin
		dbg_uart_bytes_count <= dbg_uart_bytes_count_uartwishbonebridge_next_value0;
	end
	if (dbg_uart_words_count_uartwishbonebridge_next_value_ce1) begin
		dbg_uart_words_count <= dbg_uart_words_count_uartwishbonebridge_next_value1;
	end
	if (dbg_uart_cmd_uartwishbonebridge_next_value_ce2) begin
		dbg_uart_cmd <= dbg_uart_cmd_uartwishbonebridge_next_value2;
	end
	if (dbg_uart_length_uartwishbonebridge_next_value_ce3) begin
		dbg_uart_length <= dbg_uart_length_uartwishbonebridge_next_value3;
	end
	if (dbg_uart_address_uartwishbonebridge_next_value_ce4) begin
		dbg_uart_address <= dbg_uart_address_uartwishbonebridge_next_value4;
	end
	if (dbg_uart_incr_uartwishbonebridge_next_value_ce5) begin
		dbg_uart_incr <= dbg_uart_incr_uartwishbonebridge_next_value5;
	end
	if (dbg_uart_data_uartwishbonebridge_next_value_ce6) begin
		dbg_uart_data <= dbg_uart_data_uartwishbonebridge_next_value6;
	end
	if (dbg_uart_reset) begin
		dbg_uart_incr <= 1'd0;
		uartwishbonebridge_state <= 3'd0;
	end
	if (dbg_uart_wait) begin
		if ((~dbg_uart_done)) begin
			dbg_uart_count <= (dbg_uart_count - 1'd1);
		end
	end else begin
		dbg_uart_count <= 20'd1000000;
	end
	gpioin0_gpioin0_in_pads_n_d <= gpioin0_in_status;
	if (gpioin0_gpioin0_clear) begin
		gpioin0_gpioin0_pending <= 1'd0;
	end
	gpioin0_gpioin0_trigger_d <= gpioin0_gpioin0_trigger;
	if ((gpioin0_gpioin0_trigger & (~gpioin0_gpioin0_trigger_d))) begin
		gpioin0_gpioin0_pending <= 1'd1;
	end
	gpioin1_gpioin1_in_pads_n_d <= gpioin1_in_status;
	if (gpioin1_gpioin1_clear) begin
		gpioin1_gpioin1_pending <= 1'd0;
	end
	gpioin1_gpioin1_trigger_d <= gpioin1_gpioin1_trigger;
	if ((gpioin1_gpioin1_trigger & (~gpioin1_gpioin1_trigger_d))) begin
		gpioin1_gpioin1_pending <= 1'd1;
	end
	gpioin2_gpioin2_in_pads_n_d <= gpioin2_in_status;
	if (gpioin2_gpioin2_clear) begin
		gpioin2_gpioin2_pending <= 1'd0;
	end
	gpioin2_gpioin2_trigger_d <= gpioin2_gpioin2_trigger;
	if ((gpioin2_gpioin2_trigger & (~gpioin2_gpioin2_trigger_d))) begin
		gpioin2_gpioin2_pending <= 1'd1;
	end
	gpioin3_gpioin3_in_pads_n_d <= gpioin3_in_status;
	if (gpioin3_gpioin3_clear) begin
		gpioin3_gpioin3_pending <= 1'd0;
	end
	gpioin3_gpioin3_trigger_d <= gpioin3_gpioin3_trigger;
	if ((gpioin3_gpioin3_trigger & (~gpioin3_gpioin3_trigger_d))) begin
		gpioin3_gpioin3_pending <= 1'd1;
	end
	gpioin4_gpioin4_in_pads_n_d <= gpioin4_in_status;
	if (gpioin4_gpioin4_clear) begin
		gpioin4_gpioin4_pending <= 1'd0;
	end
	gpioin4_gpioin4_trigger_d <= gpioin4_gpioin4_trigger;
	if ((gpioin4_gpioin4_trigger & (~gpioin4_gpioin4_trigger_d))) begin
		gpioin4_gpioin4_pending <= 1'd1;
	end
	gpioin5_gpioin5_in_pads_n_d <= gpioin5_in_status;
	if (gpioin5_gpioin5_clear) begin
		gpioin5_gpioin5_pending <= 1'd0;
	end
	gpioin5_gpioin5_trigger_d <= gpioin5_gpioin5_trigger;
	if ((gpioin5_gpioin5_trigger & (~gpioin5_gpioin5_trigger_d))) begin
		gpioin5_gpioin5_pending <= 1'd1;
	end
	state <= next_state;
	case (grant)
		1'd0: begin
			if ((~request[0])) begin
				if (request[1]) begin
					grant <= 1'd1;
				end else begin
					if (request[2]) begin
						grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~request[1])) begin
				if (request[2]) begin
					grant <= 2'd2;
				end else begin
					if (request[0]) begin
						grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~request[2])) begin
				if (request[0]) begin
					grant <= 1'd0;
				end else begin
					if (request[1]) begin
						grant <= 1'd1;
					end
				end
			end
		end
	endcase
	slave_sel_r <= slave_sel;
	if (wait_1) begin
		if ((~done)) begin
			count <= (count - 1'd1);
		end
	end else begin
		count <= 20'd1000000;
	end
	interface0_bank_bus_dat_r <= 1'd0;
	if (csrbank0_sel) begin
		case (interface0_bank_bus_adr[8:0])
			1'd0: begin
				interface0_bank_bus_dat_r <= csrbank0_reset0_w;
			end
			1'd1: begin
				interface0_bank_bus_dat_r <= csrbank0_scratch0_w;
			end
			2'd2: begin
				interface0_bank_bus_dat_r <= csrbank0_bus_errors_w;
			end
		endcase
	end
	if (csrbank0_reset0_re) begin
		mgmtsoc_reset_storage[1:0] <= csrbank0_reset0_r;
	end
	mgmtsoc_reset_re <= csrbank0_reset0_re;
	if (csrbank0_scratch0_re) begin
		mgmtsoc_scratch_storage[31:0] <= csrbank0_scratch0_r;
	end
	mgmtsoc_scratch_re <= csrbank0_scratch0_re;
	mgmtsoc_bus_errors_re <= csrbank0_bus_errors_re;
	interface1_bank_bus_dat_r <= 1'd0;
	if (csrbank1_sel) begin
		case (interface1_bank_bus_adr[8:0])
			1'd0: begin
				interface1_bank_bus_dat_r <= csrbank1_out0_w;
			end
		endcase
	end
	if (csrbank1_out0_re) begin
		debug_mode_storage <= csrbank1_out0_r;
	end
	debug_mode_re <= csrbank1_out0_re;
	interface2_bank_bus_dat_r <= 1'd0;
	if (csrbank2_sel) begin
		case (interface2_bank_bus_adr[8:0])
			1'd0: begin
				interface2_bank_bus_dat_r <= csrbank2_out0_w;
			end
		endcase
	end
	if (csrbank2_out0_re) begin
		debug_oeb_storage <= csrbank2_out0_r;
	end
	debug_oeb_re <= csrbank2_out0_re;
	interface3_bank_bus_dat_r <= 1'd0;
	if (csrbank3_sel) begin
		case (interface3_bank_bus_adr[8:0])
			1'd0: begin
				interface3_bank_bus_dat_r <= csrbank3_mmap_dummy_bits0_w;
			end
			1'd1: begin
				interface3_bank_bus_dat_r <= csrbank3_master_cs0_w;
			end
			2'd2: begin
				interface3_bank_bus_dat_r <= csrbank3_master_phyconfig0_w;
			end
			2'd3: begin
				interface3_bank_bus_dat_r <= mgmtsoc_master_rxtx_w;
			end
			3'd4: begin
				interface3_bank_bus_dat_r <= csrbank3_master_status_w;
			end
		endcase
	end
	if (csrbank3_mmap_dummy_bits0_re) begin
		mgmtsoc_litespimmap_storage[7:0] <= csrbank3_mmap_dummy_bits0_r;
	end
	mgmtsoc_litespimmap_re <= csrbank3_mmap_dummy_bits0_re;
	if (csrbank3_master_cs0_re) begin
		mgmtsoc_master_cs_storage <= csrbank3_master_cs0_r;
	end
	mgmtsoc_master_cs_re <= csrbank3_master_cs0_re;
	if (csrbank3_master_phyconfig0_re) begin
		mgmtsoc_master_phyconfig_storage[23:0] <= csrbank3_master_phyconfig0_r;
	end
	mgmtsoc_master_phyconfig_re <= csrbank3_master_phyconfig0_re;
	mgmtsoc_master_status_re <= csrbank3_master_status_re;
	interface4_bank_bus_dat_r <= 1'd0;
	if (csrbank4_sel) begin
		case (interface4_bank_bus_adr[8:0])
			1'd0: begin
				interface4_bank_bus_dat_r <= csrbank4_clk_divisor0_w;
			end
		endcase
	end
	if (csrbank4_clk_divisor0_re) begin
		mgmtsoc_litespisdrphycore_storage[7:0] <= csrbank4_clk_divisor0_r;
	end
	mgmtsoc_litespisdrphycore_re <= csrbank4_clk_divisor0_re;
	interface5_bank_bus_dat_r <= 1'd0;
	if (csrbank5_sel) begin
		case (interface5_bank_bus_adr[8:0])
			1'd0: begin
				interface5_bank_bus_dat_r <= csrbank5_mode10_w;
			end
			1'd1: begin
				interface5_bank_bus_dat_r <= csrbank5_mode00_w;
			end
			2'd2: begin
				interface5_bank_bus_dat_r <= csrbank5_ien0_w;
			end
			2'd3: begin
				interface5_bank_bus_dat_r <= csrbank5_oe0_w;
			end
			3'd4: begin
				interface5_bank_bus_dat_r <= csrbank5_in_w;
			end
			3'd5: begin
				interface5_bank_bus_dat_r <= csrbank5_out0_w;
			end
		endcase
	end
	if (csrbank5_mode10_re) begin
		gpio_mode1_storage <= csrbank5_mode10_r;
	end
	gpio_mode1_re <= csrbank5_mode10_re;
	if (csrbank5_mode00_re) begin
		gpio_mode0_storage <= csrbank5_mode00_r;
	end
	gpio_mode0_re <= csrbank5_mode00_re;
	if (csrbank5_ien0_re) begin
		gpio_ien_storage <= csrbank5_ien0_r;
	end
	gpio_ien_re <= csrbank5_ien0_re;
	if (csrbank5_oe0_re) begin
		gpio_oe_storage <= csrbank5_oe0_r;
	end
	gpio_oe_re <= csrbank5_oe0_re;
	gpio_in_re <= csrbank5_in_re;
	if (csrbank5_out0_re) begin
		gpio_out_storage <= csrbank5_out0_r;
	end
	gpio_out_re <= csrbank5_out0_re;
	interface6_bank_bus_dat_r <= 1'd0;
	if (csrbank6_sel) begin
		case (interface6_bank_bus_adr[8:0])
			1'd0: begin
				interface6_bank_bus_dat_r <= csrbank6_ien3_w;
			end
			1'd1: begin
				interface6_bank_bus_dat_r <= csrbank6_ien2_w;
			end
			2'd2: begin
				interface6_bank_bus_dat_r <= csrbank6_ien1_w;
			end
			2'd3: begin
				interface6_bank_bus_dat_r <= csrbank6_ien0_w;
			end
			3'd4: begin
				interface6_bank_bus_dat_r <= csrbank6_oe3_w;
			end
			3'd5: begin
				interface6_bank_bus_dat_r <= csrbank6_oe2_w;
			end
			3'd6: begin
				interface6_bank_bus_dat_r <= csrbank6_oe1_w;
			end
			3'd7: begin
				interface6_bank_bus_dat_r <= csrbank6_oe0_w;
			end
			4'd8: begin
				interface6_bank_bus_dat_r <= csrbank6_in3_w;
			end
			4'd9: begin
				interface6_bank_bus_dat_r <= csrbank6_in2_w;
			end
			4'd10: begin
				interface6_bank_bus_dat_r <= csrbank6_in1_w;
			end
			4'd11: begin
				interface6_bank_bus_dat_r <= csrbank6_in0_w;
			end
			4'd12: begin
				interface6_bank_bus_dat_r <= csrbank6_out3_w;
			end
			4'd13: begin
				interface6_bank_bus_dat_r <= csrbank6_out2_w;
			end
			4'd14: begin
				interface6_bank_bus_dat_r <= csrbank6_out1_w;
			end
			4'd15: begin
				interface6_bank_bus_dat_r <= csrbank6_out0_w;
			end
		endcase
	end
	if (csrbank6_ien3_re) begin
		la_ien_storage[127:96] <= csrbank6_ien3_r;
	end
	if (csrbank6_ien2_re) begin
		la_ien_storage[95:64] <= csrbank6_ien2_r;
	end
	if (csrbank6_ien1_re) begin
		la_ien_storage[63:32] <= csrbank6_ien1_r;
	end
	if (csrbank6_ien0_re) begin
		la_ien_storage[31:0] <= csrbank6_ien0_r;
	end
	la_ien_re <= csrbank6_ien0_re;
	if (csrbank6_oe3_re) begin
		la_oe_storage[127:96] <= csrbank6_oe3_r;
	end
	if (csrbank6_oe2_re) begin
		la_oe_storage[95:64] <= csrbank6_oe2_r;
	end
	if (csrbank6_oe1_re) begin
		la_oe_storage[63:32] <= csrbank6_oe1_r;
	end
	if (csrbank6_oe0_re) begin
		la_oe_storage[31:0] <= csrbank6_oe0_r;
	end
	la_oe_re <= csrbank6_oe0_re;
	la_in_re <= csrbank6_in0_re;
	if (csrbank6_out3_re) begin
		la_out_storage[127:96] <= csrbank6_out3_r;
	end
	if (csrbank6_out2_re) begin
		la_out_storage[95:64] <= csrbank6_out2_r;
	end
	if (csrbank6_out1_re) begin
		la_out_storage[63:32] <= csrbank6_out1_r;
	end
	if (csrbank6_out0_re) begin
		la_out_storage[31:0] <= csrbank6_out0_r;
	end
	la_out_re <= csrbank6_out0_re;
	interface7_bank_bus_dat_r <= 1'd0;
	if (csrbank7_sel) begin
		case (interface7_bank_bus_adr[8:0])
			1'd0: begin
				interface7_bank_bus_dat_r <= csrbank7_out0_w;
			end
		endcase
	end
	if (csrbank7_out0_re) begin
		mprj_wb_iena_storage <= csrbank7_out0_r;
	end
	mprj_wb_iena_re <= csrbank7_out0_re;
	interface8_bank_bus_dat_r <= 1'd0;
	if (csrbank8_sel) begin
		case (interface8_bank_bus_adr[8:0])
			1'd0: begin
				interface8_bank_bus_dat_r <= csrbank8_out0_w;
			end
		endcase
	end
	if (csrbank8_out0_re) begin
		spi_enabled_storage <= csrbank8_out0_r;
	end
	spi_enabled_re <= csrbank8_out0_re;
	interface9_bank_bus_dat_r <= 1'd0;
	if (csrbank9_sel) begin
		case (interface9_bank_bus_adr[8:0])
			1'd0: begin
				interface9_bank_bus_dat_r <= csrbank9_control0_w;
			end
			1'd1: begin
				interface9_bank_bus_dat_r <= csrbank9_status_w;
			end
			2'd2: begin
				interface9_bank_bus_dat_r <= csrbank9_mosi0_w;
			end
			2'd3: begin
				interface9_bank_bus_dat_r <= csrbank9_miso_w;
			end
			3'd4: begin
				interface9_bank_bus_dat_r <= csrbank9_cs0_w;
			end
			3'd5: begin
				interface9_bank_bus_dat_r <= csrbank9_loopback0_w;
			end
			3'd6: begin
				interface9_bank_bus_dat_r <= csrbank9_clk_divider0_w;
			end
		endcase
	end
	if (csrbank9_control0_re) begin
		spi_master_control_storage[15:0] <= csrbank9_control0_r;
	end
	spi_master_control_re <= csrbank9_control0_re;
	spi_master_status_re <= csrbank9_status_re;
	if (csrbank9_mosi0_re) begin
		spi_master_mosi_storage[7:0] <= csrbank9_mosi0_r;
	end
	spi_master_mosi_re <= csrbank9_mosi0_re;
	spi_master_miso_re <= csrbank9_miso_re;
	if (csrbank9_cs0_re) begin
		spi_master_cs_storage[16:0] <= csrbank9_cs0_r;
	end
	spi_master_cs_re <= csrbank9_cs0_re;
	if (csrbank9_loopback0_re) begin
		spi_master_loopback_storage <= csrbank9_loopback0_r;
	end
	spi_master_loopback_re <= csrbank9_loopback0_re;
	if (csrbank9_clk_divider0_re) begin
		spimaster_storage[15:0] <= csrbank9_clk_divider0_r;
	end
	spimaster_re <= csrbank9_clk_divider0_re;
	interface10_bank_bus_dat_r <= 1'd0;
	if (csrbank10_sel) begin
		case (interface10_bank_bus_adr[8:0])
			1'd0: begin
				interface10_bank_bus_dat_r <= csrbank10_load0_w;
			end
			1'd1: begin
				interface10_bank_bus_dat_r <= csrbank10_reload0_w;
			end
			2'd2: begin
				interface10_bank_bus_dat_r <= csrbank10_en0_w;
			end
			2'd3: begin
				interface10_bank_bus_dat_r <= csrbank10_update_value0_w;
			end
			3'd4: begin
				interface10_bank_bus_dat_r <= csrbank10_value_w;
			end
			3'd5: begin
				interface10_bank_bus_dat_r <= csrbank10_ev_status_w;
			end
			3'd6: begin
				interface10_bank_bus_dat_r <= csrbank10_ev_pending_w;
			end
			3'd7: begin
				interface10_bank_bus_dat_r <= csrbank10_ev_enable0_w;
			end
		endcase
	end
	if (csrbank10_load0_re) begin
		mgmtsoc_load_storage[31:0] <= csrbank10_load0_r;
	end
	mgmtsoc_load_re <= csrbank10_load0_re;
	if (csrbank10_reload0_re) begin
		mgmtsoc_reload_storage[31:0] <= csrbank10_reload0_r;
	end
	mgmtsoc_reload_re <= csrbank10_reload0_re;
	if (csrbank10_en0_re) begin
		mgmtsoc_en_storage <= csrbank10_en0_r;
	end
	mgmtsoc_en_re <= csrbank10_en0_re;
	if (csrbank10_update_value0_re) begin
		mgmtsoc_update_value_storage <= csrbank10_update_value0_r;
	end
	mgmtsoc_update_value_re <= csrbank10_update_value0_re;
	mgmtsoc_value_re <= csrbank10_value_re;
	mgmtsoc_status_re <= csrbank10_ev_status_re;
	if (csrbank10_ev_pending_re) begin
		mgmtsoc_pending_r <= csrbank10_ev_pending_r;
	end
	mgmtsoc_pending_re <= csrbank10_ev_pending_re;
	if (csrbank10_ev_enable0_re) begin
		mgmtsoc_enable_storage <= csrbank10_ev_enable0_r;
	end
	mgmtsoc_enable_re <= csrbank10_ev_enable0_re;
	interface11_bank_bus_dat_r <= 1'd0;
	if (csrbank11_sel) begin
		case (interface11_bank_bus_adr[8:0])
			1'd0: begin
				interface11_bank_bus_dat_r <= uart_rxtx_w;
			end
			1'd1: begin
				interface11_bank_bus_dat_r <= csrbank11_txfull_w;
			end
			2'd2: begin
				interface11_bank_bus_dat_r <= csrbank11_rxempty_w;
			end
			2'd3: begin
				interface11_bank_bus_dat_r <= csrbank11_ev_status_w;
			end
			3'd4: begin
				interface11_bank_bus_dat_r <= csrbank11_ev_pending_w;
			end
			3'd5: begin
				interface11_bank_bus_dat_r <= csrbank11_ev_enable0_w;
			end
			3'd6: begin
				interface11_bank_bus_dat_r <= csrbank11_txempty_w;
			end
			3'd7: begin
				interface11_bank_bus_dat_r <= csrbank11_rxfull_w;
			end
		endcase
	end
	uart_txfull_re <= csrbank11_txfull_re;
	uart_rxempty_re <= csrbank11_rxempty_re;
	uart_status_re <= csrbank11_ev_status_re;
	if (csrbank11_ev_pending_re) begin
		uart_pending_r[1:0] <= csrbank11_ev_pending_r;
	end
	uart_pending_re <= csrbank11_ev_pending_re;
	if (csrbank11_ev_enable0_re) begin
		uart_enable_storage[1:0] <= csrbank11_ev_enable0_r;
	end
	uart_enable_re <= csrbank11_ev_enable0_re;
	uart_txempty_re <= csrbank11_txempty_re;
	uart_rxfull_re <= csrbank11_rxfull_re;
	interface12_bank_bus_dat_r <= 1'd0;
	if (csrbank12_sel) begin
		case (interface12_bank_bus_adr[8:0])
			1'd0: begin
				interface12_bank_bus_dat_r <= csrbank12_out0_w;
			end
		endcase
	end
	if (csrbank12_out0_re) begin
		uart_enabled_storage <= csrbank12_out0_r;
	end
	uart_enabled_re <= csrbank12_out0_re;
	interface13_bank_bus_dat_r <= 1'd0;
	if (csrbank13_sel) begin
		case (interface13_bank_bus_adr[8:0])
			1'd0: begin
				interface13_bank_bus_dat_r <= csrbank13_in_w;
			end
			1'd1: begin
				interface13_bank_bus_dat_r <= csrbank13_mode0_w;
			end
			2'd2: begin
				interface13_bank_bus_dat_r <= csrbank13_edge0_w;
			end
			2'd3: begin
				interface13_bank_bus_dat_r <= csrbank13_ev_status_w;
			end
			3'd4: begin
				interface13_bank_bus_dat_r <= csrbank13_ev_pending_w;
			end
			3'd5: begin
				interface13_bank_bus_dat_r <= csrbank13_ev_enable0_w;
			end
		endcase
	end
	gpioin0_in_re <= csrbank13_in_re;
	if (csrbank13_mode0_re) begin
		gpioin0_gpioin0_mode_storage <= csrbank13_mode0_r;
	end
	gpioin0_gpioin0_mode_re <= csrbank13_mode0_re;
	if (csrbank13_edge0_re) begin
		gpioin0_gpioin0_edge_storage <= csrbank13_edge0_r;
	end
	gpioin0_gpioin0_edge_re <= csrbank13_edge0_re;
	gpioin0_status_re <= csrbank13_ev_status_re;
	if (csrbank13_ev_pending_re) begin
		gpioin0_pending_r <= csrbank13_ev_pending_r;
	end
	gpioin0_pending_re <= csrbank13_ev_pending_re;
	if (csrbank13_ev_enable0_re) begin
		gpioin0_enable_storage <= csrbank13_ev_enable0_r;
	end
	gpioin0_enable_re <= csrbank13_ev_enable0_re;
	interface14_bank_bus_dat_r <= 1'd0;
	if (csrbank14_sel) begin
		case (interface14_bank_bus_adr[8:0])
			1'd0: begin
				interface14_bank_bus_dat_r <= csrbank14_in_w;
			end
			1'd1: begin
				interface14_bank_bus_dat_r <= csrbank14_mode0_w;
			end
			2'd2: begin
				interface14_bank_bus_dat_r <= csrbank14_edge0_w;
			end
			2'd3: begin
				interface14_bank_bus_dat_r <= csrbank14_ev_status_w;
			end
			3'd4: begin
				interface14_bank_bus_dat_r <= csrbank14_ev_pending_w;
			end
			3'd5: begin
				interface14_bank_bus_dat_r <= csrbank14_ev_enable0_w;
			end
		endcase
	end
	gpioin1_in_re <= csrbank14_in_re;
	if (csrbank14_mode0_re) begin
		gpioin1_gpioin1_mode_storage <= csrbank14_mode0_r;
	end
	gpioin1_gpioin1_mode_re <= csrbank14_mode0_re;
	if (csrbank14_edge0_re) begin
		gpioin1_gpioin1_edge_storage <= csrbank14_edge0_r;
	end
	gpioin1_gpioin1_edge_re <= csrbank14_edge0_re;
	gpioin1_status_re <= csrbank14_ev_status_re;
	if (csrbank14_ev_pending_re) begin
		gpioin1_pending_r <= csrbank14_ev_pending_r;
	end
	gpioin1_pending_re <= csrbank14_ev_pending_re;
	if (csrbank14_ev_enable0_re) begin
		gpioin1_enable_storage <= csrbank14_ev_enable0_r;
	end
	gpioin1_enable_re <= csrbank14_ev_enable0_re;
	interface15_bank_bus_dat_r <= 1'd0;
	if (csrbank15_sel) begin
		case (interface15_bank_bus_adr[8:0])
			1'd0: begin
				interface15_bank_bus_dat_r <= csrbank15_in_w;
			end
			1'd1: begin
				interface15_bank_bus_dat_r <= csrbank15_mode0_w;
			end
			2'd2: begin
				interface15_bank_bus_dat_r <= csrbank15_edge0_w;
			end
			2'd3: begin
				interface15_bank_bus_dat_r <= csrbank15_ev_status_w;
			end
			3'd4: begin
				interface15_bank_bus_dat_r <= csrbank15_ev_pending_w;
			end
			3'd5: begin
				interface15_bank_bus_dat_r <= csrbank15_ev_enable0_w;
			end
		endcase
	end
	gpioin2_in_re <= csrbank15_in_re;
	if (csrbank15_mode0_re) begin
		gpioin2_gpioin2_mode_storage <= csrbank15_mode0_r;
	end
	gpioin2_gpioin2_mode_re <= csrbank15_mode0_re;
	if (csrbank15_edge0_re) begin
		gpioin2_gpioin2_edge_storage <= csrbank15_edge0_r;
	end
	gpioin2_gpioin2_edge_re <= csrbank15_edge0_re;
	gpioin2_status_re <= csrbank15_ev_status_re;
	if (csrbank15_ev_pending_re) begin
		gpioin2_pending_r <= csrbank15_ev_pending_r;
	end
	gpioin2_pending_re <= csrbank15_ev_pending_re;
	if (csrbank15_ev_enable0_re) begin
		gpioin2_enable_storage <= csrbank15_ev_enable0_r;
	end
	gpioin2_enable_re <= csrbank15_ev_enable0_re;
	interface16_bank_bus_dat_r <= 1'd0;
	if (csrbank16_sel) begin
		case (interface16_bank_bus_adr[8:0])
			1'd0: begin
				interface16_bank_bus_dat_r <= csrbank16_in_w;
			end
			1'd1: begin
				interface16_bank_bus_dat_r <= csrbank16_mode0_w;
			end
			2'd2: begin
				interface16_bank_bus_dat_r <= csrbank16_edge0_w;
			end
			2'd3: begin
				interface16_bank_bus_dat_r <= csrbank16_ev_status_w;
			end
			3'd4: begin
				interface16_bank_bus_dat_r <= csrbank16_ev_pending_w;
			end
			3'd5: begin
				interface16_bank_bus_dat_r <= csrbank16_ev_enable0_w;
			end
		endcase
	end
	gpioin3_in_re <= csrbank16_in_re;
	if (csrbank16_mode0_re) begin
		gpioin3_gpioin3_mode_storage <= csrbank16_mode0_r;
	end
	gpioin3_gpioin3_mode_re <= csrbank16_mode0_re;
	if (csrbank16_edge0_re) begin
		gpioin3_gpioin3_edge_storage <= csrbank16_edge0_r;
	end
	gpioin3_gpioin3_edge_re <= csrbank16_edge0_re;
	gpioin3_status_re <= csrbank16_ev_status_re;
	if (csrbank16_ev_pending_re) begin
		gpioin3_pending_r <= csrbank16_ev_pending_r;
	end
	gpioin3_pending_re <= csrbank16_ev_pending_re;
	if (csrbank16_ev_enable0_re) begin
		gpioin3_enable_storage <= csrbank16_ev_enable0_r;
	end
	gpioin3_enable_re <= csrbank16_ev_enable0_re;
	interface17_bank_bus_dat_r <= 1'd0;
	if (csrbank17_sel) begin
		case (interface17_bank_bus_adr[8:0])
			1'd0: begin
				interface17_bank_bus_dat_r <= csrbank17_in_w;
			end
			1'd1: begin
				interface17_bank_bus_dat_r <= csrbank17_mode0_w;
			end
			2'd2: begin
				interface17_bank_bus_dat_r <= csrbank17_edge0_w;
			end
			2'd3: begin
				interface17_bank_bus_dat_r <= csrbank17_ev_status_w;
			end
			3'd4: begin
				interface17_bank_bus_dat_r <= csrbank17_ev_pending_w;
			end
			3'd5: begin
				interface17_bank_bus_dat_r <= csrbank17_ev_enable0_w;
			end
		endcase
	end
	gpioin4_in_re <= csrbank17_in_re;
	if (csrbank17_mode0_re) begin
		gpioin4_gpioin4_mode_storage <= csrbank17_mode0_r;
	end
	gpioin4_gpioin4_mode_re <= csrbank17_mode0_re;
	if (csrbank17_edge0_re) begin
		gpioin4_gpioin4_edge_storage <= csrbank17_edge0_r;
	end
	gpioin4_gpioin4_edge_re <= csrbank17_edge0_re;
	gpioin4_status_re <= csrbank17_ev_status_re;
	if (csrbank17_ev_pending_re) begin
		gpioin4_pending_r <= csrbank17_ev_pending_r;
	end
	gpioin4_pending_re <= csrbank17_ev_pending_re;
	if (csrbank17_ev_enable0_re) begin
		gpioin4_enable_storage <= csrbank17_ev_enable0_r;
	end
	gpioin4_enable_re <= csrbank17_ev_enable0_re;
	interface18_bank_bus_dat_r <= 1'd0;
	if (csrbank18_sel) begin
		case (interface18_bank_bus_adr[8:0])
			1'd0: begin
				interface18_bank_bus_dat_r <= csrbank18_in_w;
			end
			1'd1: begin
				interface18_bank_bus_dat_r <= csrbank18_mode0_w;
			end
			2'd2: begin
				interface18_bank_bus_dat_r <= csrbank18_edge0_w;
			end
			2'd3: begin
				interface18_bank_bus_dat_r <= csrbank18_ev_status_w;
			end
			3'd4: begin
				interface18_bank_bus_dat_r <= csrbank18_ev_pending_w;
			end
			3'd5: begin
				interface18_bank_bus_dat_r <= csrbank18_ev_enable0_w;
			end
		endcase
	end
	gpioin5_in_re <= csrbank18_in_re;
	if (csrbank18_mode0_re) begin
		gpioin5_gpioin5_mode_storage <= csrbank18_mode0_r;
	end
	gpioin5_gpioin5_mode_re <= csrbank18_mode0_re;
	if (csrbank18_edge0_re) begin
		gpioin5_gpioin5_edge_storage <= csrbank18_edge0_r;
	end
	gpioin5_gpioin5_edge_re <= csrbank18_edge0_re;
	gpioin5_status_re <= csrbank18_ev_status_re;
	if (csrbank18_ev_pending_re) begin
		gpioin5_pending_r <= csrbank18_ev_pending_r;
	end
	gpioin5_pending_re <= csrbank18_ev_pending_re;
	if (csrbank18_ev_enable0_re) begin
		gpioin5_enable_storage <= csrbank18_ev_enable0_r;
	end
	gpioin5_enable_re <= csrbank18_ev_enable0_re;
	interface19_bank_bus_dat_r <= 1'd0;
	if (csrbank19_sel) begin
		case (interface19_bank_bus_adr[8:0])
			1'd0: begin
				interface19_bank_bus_dat_r <= csrbank19_out0_w;
			end
		endcase
	end
	if (csrbank19_out0_re) begin
		user_irq_ena_storage[2:0] <= csrbank19_out0_r;
	end
	user_irq_ena_re <= csrbank19_out0_re;
	if (sys_rst) begin
	    // ****** added to correct GL testbench failure
        dbg_uart_tx_data <= 8'd0;
        dbg_uart_tx_count <= 4'd0;
        dbg_uart_tx_tick <= 1'd0;
        dbg_uart_tx_phase <= 32'd0;
        dbg_uart_rx_tick <= 1'd0;
        dbg_uart_rx_phase <= 32'd0;
        dbg_uart_rx_rx_d <= 1'd0;
        dbg_uart_cmd <= 8'd0;
        dbg_uart_incr <= 1'd0;
        dbg_uart_address <= 32'd0;
        dbg_uart_data <= 32'd0;
        dbg_uart_bytes_count <= 2'd0;
        dbg_uart_words_count <= 8'd0;
        dbg_uart_count <= 20'd1000000;
	    // ******
		mgmtsoc_reset_storage <= 2'd0;
		mgmtsoc_reset_re <= 1'd0;
		mgmtsoc_scratch_storage <= 32'd305419896;
		mgmtsoc_scratch_re <= 1'd0;
		mgmtsoc_bus_errors_re <= 1'd0;
		mgmtsoc_bus_errors <= 32'd0;
		mgmtsoc_vexriscv_debug_reset <= 1'd0;
		mgmtsoc_vexriscv_ibus_err <= 1'd0;
		mgmtsoc_vexriscv_dbus_err <= 1'd0;
		mgmtsoc_vexriscv_i_cmd_valid <= 1'd0;
		mgmtsoc_vexriscv_i_cmd_payload_wr <= 1'd0;
		mgmtsoc_vexriscv_i_cmd_payload_address <= 8'd0;
		mgmtsoc_vexriscv_i_cmd_payload_data <= 32'd0;
		mgmtsoc_vexriscv_reset_debug_logic <= 1'd0;
		mgmtsoc_vexriscv_transfer_complete <= 1'd0;
		mgmtsoc_vexriscv_transfer_in_progress <= 1'd0;
		mgmtsoc_vexriscv_transfer_wait_for_ack <= 1'd0;
		mgmtsoc_vexriscv_debug_bus_ack <= 1'd0;
		mgmtsoc_load_storage <= 32'd0;
		mgmtsoc_load_re <= 1'd0;
		mgmtsoc_reload_storage <= 32'd0;
		mgmtsoc_reload_re <= 1'd0;
		mgmtsoc_en_storage <= 1'd0;
		mgmtsoc_en_re <= 1'd0;
		mgmtsoc_update_value_storage <= 1'd0;
		mgmtsoc_update_value_re <= 1'd0;
		mgmtsoc_value_status <= 32'd0;
		mgmtsoc_value_re <= 1'd0;
		mgmtsoc_zero_pending <= 1'd0;
		mgmtsoc_zero_trigger_d <= 1'd0;
		mgmtsoc_status_re <= 1'd0;
		mgmtsoc_pending_re <= 1'd0;
		mgmtsoc_pending_r <= 1'd0;
		mgmtsoc_enable_storage <= 1'd0;
		mgmtsoc_enable_re <= 1'd0;
		mgmtsoc_value <= 32'd0;
		dff_bus_ack <= 1'd0;
		dff2_bus_ack <= 1'd0;
		mgmtsoc_litespisdrphycore_storage <= 8'd1;
		mgmtsoc_litespisdrphycore_re <= 1'd0;
		mgmtsoc_litespisdrphycore_cnt <= 8'd0;
		mgmtsoc_litespisdrphycore_clk <= 1'd0;
		mgmtsoc_litespisdrphycore_posedge_reg <= 1'd0;
		mgmtsoc_litespisdrphycore_posedge_reg2 <= 1'd0;
		mgmtsoc_litespisdrphycore_count <= 4'd11;
		mgmtsoc_litespimmap_burst_cs <= 1'd0;
		mgmtsoc_litespimmap_count <= 9'd256;
		mgmtsoc_litespimmap_storage <= 8'd0;
		mgmtsoc_litespimmap_re <= 1'd0;
		mgmtsoc_master_cs_storage <= 1'd0;
		mgmtsoc_master_cs_re <= 1'd0;
		mgmtsoc_master_phyconfig_storage <= 24'd0;
		mgmtsoc_master_phyconfig_re <= 1'd0;
		mgmtsoc_master_status_re <= 1'd0;
		mgmtsoc_master_tx_fifo_source_valid <= 1'd0;
		mgmtsoc_master_tx_fifo_source_payload_data <= 32'd0;
		mgmtsoc_master_tx_fifo_source_payload_len <= 6'd0;
		mgmtsoc_master_tx_fifo_source_payload_width <= 4'd0;
		mgmtsoc_master_tx_fifo_source_payload_mask <= 8'd0;
		mgmtsoc_master_rx_fifo_source_valid <= 1'd0;
		mgmtsoc_master_rx_fifo_source_payload_data <= 32'd0;
		spi_clk <= 1'd0;
		spi_cs_n <= 1'd0;
		spi_mosi <= 1'd0;
		spi_master_miso <= 8'd0;
		spi_master_control_storage <= 16'd0;
		spi_master_control_re <= 1'd0;
		spi_master_status_re <= 1'd0;
		spi_master_mosi_re <= 1'd0;
		spi_master_miso_re <= 1'd0;
		spi_master_cs_storage <= 17'd1;
		spi_master_cs_re <= 1'd0;
		spi_master_loopback_storage <= 1'd0;
		spi_master_loopback_re <= 1'd0;
		spi_master_count <= 3'd0;
		spi_master_clk_divider1 <= 16'd0;
		spi_master_mosi_data <= 8'd0;
		spi_master_mosi_sel <= 3'd0;
		spi_master_miso_data <= 8'd0;
		spimaster_storage <= 16'd100;
		spimaster_re <= 1'd0;
		mprj_wb_iena_storage <= 1'd0;
		mprj_wb_iena_re <= 1'd0;
		sys_uart_tx <= 1'd1;
		uart_phy_tx_tick <= 1'd0;
		uart_phy_rx_tick <= 1'd0;
		uart_phy_rx_rx_d <= 1'd0;
		uart_txfull_re <= 1'd0;
		uart_rxempty_re <= 1'd0;
		uart_tx_pending <= 1'd0;
		uart_tx_trigger_d <= 1'd0;
		uart_rx_pending <= 1'd0;
		uart_rx_trigger_d <= 1'd0;
		uart_status_re <= 1'd0;
		uart_pending_re <= 1'd0;
		uart_pending_r <= 2'd0;
		uart_enable_storage <= 2'd0;
		uart_enable_re <= 1'd0;
		uart_txempty_re <= 1'd0;
		uart_rxfull_re <= 1'd0;
		uart_tx_fifo_readable <= 1'd0;
		uart_tx_fifo_level0 <= 5'd0;
		uart_tx_fifo_produce <= 4'd0;
		uart_tx_fifo_consume <= 4'd0;
		uart_rx_fifo_readable <= 1'd0;
		uart_rx_fifo_level0 <= 5'd0;
		uart_rx_fifo_produce <= 4'd0;
		uart_rx_fifo_consume <= 4'd0;
		dbg_uart_dbg_uart_tx <= 1'd1;
		dbg_uart_tx_tick <= 1'd0;
		dbg_uart_rx_tick <= 1'd0;
		dbg_uart_rx_rx_d <= 1'd0;
		dbg_uart_incr <= 1'd0;
		dbg_uart_count <= 20'd1000000;
		debug_oeb_storage <= 1'd0;
		debug_oeb_re <= 1'd0;
		debug_mode_storage <= 1'd0;
		debug_mode_re <= 1'd0;
		uart_enabled_storage <= 1'd0;
		uart_enabled_re <= 1'd0;
		gpio_mode1_storage <= 1'd0;
		gpio_mode1_re <= 1'd0;
		gpio_mode0_storage <= 1'd0;
		gpio_mode0_re <= 1'd0;
		gpio_ien_storage <= 1'd0;
		gpio_ien_re <= 1'd0;
		gpio_oe_storage <= 1'd0;
		gpio_oe_re <= 1'd0;
		gpio_in_re <= 1'd0;
		gpio_out_storage <= 1'd0;
		gpio_out_re <= 1'd0;
		la_ien_storage <= 128'd0;
		la_ien_re <= 1'd0;
		la_oe_storage <= 128'd0;
		la_oe_re <= 1'd0;
		la_in_re <= 1'd0;
		la_out_storage <= 128'd0;
		la_out_re <= 1'd0;
		spi_enabled_storage <= 1'd0;
		spi_enabled_re <= 1'd0;
		user_irq_ena_storage <= 3'd0;
		user_irq_ena_re <= 1'd0;
		gpioin0_in_re <= 1'd0;
		gpioin0_gpioin0_mode_storage <= 1'd0;
		gpioin0_gpioin0_mode_re <= 1'd0;
		gpioin0_gpioin0_edge_storage <= 1'd0;
		gpioin0_gpioin0_edge_re <= 1'd0;
		gpioin0_gpioin0_in_pads_n_d <= 1'd0;
		gpioin0_gpioin0_pending <= 1'd0;
		gpioin0_gpioin0_trigger_d <= 1'd0;
		gpioin1_in_re <= 1'd0;
		gpioin1_gpioin1_mode_storage <= 1'd0;
		gpioin1_gpioin1_mode_re <= 1'd0;
		gpioin1_gpioin1_edge_storage <= 1'd0;
		gpioin1_gpioin1_edge_re <= 1'd0;
		gpioin1_gpioin1_in_pads_n_d <= 1'd0;
		gpioin1_gpioin1_pending <= 1'd0;
		gpioin1_gpioin1_trigger_d <= 1'd0;
		gpioin2_in_re <= 1'd0;
		gpioin2_gpioin2_mode_storage <= 1'd0;
		gpioin2_gpioin2_mode_re <= 1'd0;
		gpioin2_gpioin2_edge_storage <= 1'd0;
		gpioin2_gpioin2_edge_re <= 1'd0;
		gpioin2_gpioin2_in_pads_n_d <= 1'd0;
		gpioin2_gpioin2_pending <= 1'd0;
		gpioin2_gpioin2_trigger_d <= 1'd0;
		gpioin3_in_re <= 1'd0;
		gpioin3_gpioin3_mode_storage <= 1'd0;
		gpioin3_gpioin3_mode_re <= 1'd0;
		gpioin3_gpioin3_edge_storage <= 1'd0;
		gpioin3_gpioin3_edge_re <= 1'd0;
		gpioin3_gpioin3_in_pads_n_d <= 1'd0;
		gpioin3_gpioin3_pending <= 1'd0;
		gpioin3_gpioin3_trigger_d <= 1'd0;
		gpioin4_in_re <= 1'd0;
		gpioin4_gpioin4_mode_storage <= 1'd0;
		gpioin4_gpioin4_mode_re <= 1'd0;
		gpioin4_gpioin4_edge_storage <= 1'd0;
		gpioin4_gpioin4_edge_re <= 1'd0;
		gpioin4_gpioin4_in_pads_n_d <= 1'd0;
		gpioin4_gpioin4_pending <= 1'd0;
		gpioin4_gpioin4_trigger_d <= 1'd0;
		gpioin5_in_re <= 1'd0;
		gpioin5_gpioin5_mode_storage <= 1'd0;
		gpioin5_gpioin5_mode_re <= 1'd0;
		gpioin5_gpioin5_edge_storage <= 1'd0;
		gpioin5_gpioin5_edge_re <= 1'd0;
		gpioin5_gpioin5_in_pads_n_d <= 1'd0;
		gpioin5_gpioin5_pending <= 1'd0;
		gpioin5_gpioin5_trigger_d <= 1'd0;
		litespiphy_state <= 2'd0;
		litespi_grant <= 1'd0;
		litespi_state <= 4'd0;
		spimaster_state <= 2'd0;
		rs232phy_rs232phytx_state <= 1'd0;
		rs232phy_rs232phyrx_state <= 1'd0;
		uartwishbonebridge_rs232phytx_state <= 1'd0;
		uartwishbonebridge_rs232phyrx_state <= 1'd0;
		uartwishbonebridge_state <= 3'd0;
		gpioin0_status_re <= 1'd0;
		gpioin0_pending_re <= 1'd0;
		gpioin0_pending_r <= 1'd0;
		gpioin0_enable_storage <= 1'd0;
		gpioin0_enable_re <= 1'd0;
		gpioin1_status_re <= 1'd0;
		gpioin1_pending_re <= 1'd0;
		gpioin1_pending_r <= 1'd0;
		gpioin1_enable_storage <= 1'd0;
		gpioin1_enable_re <= 1'd0;
		gpioin2_status_re <= 1'd0;
		gpioin2_pending_re <= 1'd0;
		gpioin2_pending_r <= 1'd0;
		gpioin2_enable_storage <= 1'd0;
		gpioin2_enable_re <= 1'd0;
		gpioin3_status_re <= 1'd0;
		gpioin3_pending_re <= 1'd0;
		gpioin3_pending_r <= 1'd0;
		gpioin3_enable_storage <= 1'd0;
		gpioin3_enable_re <= 1'd0;
		gpioin4_status_re <= 1'd0;
		gpioin4_pending_re <= 1'd0;
		gpioin4_pending_r <= 1'd0;
		gpioin4_enable_storage <= 1'd0;
		gpioin4_enable_re <= 1'd0;
		gpioin5_status_re <= 1'd0;
		gpioin5_pending_re <= 1'd0;
		gpioin5_pending_r <= 1'd0;
		gpioin5_enable_storage <= 1'd0;
		gpioin5_enable_re <= 1'd0;
		grant <= 2'd0;
		slave_sel_r <= 7'd0;
		count <= 20'd1000000;
		state <= 1'd0;
	end
	multiregimpl0_regs0 <= sys_uart_rx;
	multiregimpl0_regs1 <= multiregimpl0_regs0;
	multiregimpl1_regs0 <= dbg_uart_dbg_uart_rx;
	multiregimpl1_regs1 <= multiregimpl1_regs0;
	multiregimpl2_regs0 <= gpio_in_pad;
	multiregimpl2_regs1 <= multiregimpl2_regs0;
	multiregimpl3_regs0 <= la_input[0];
	multiregimpl3_regs1 <= multiregimpl3_regs0;
	multiregimpl4_regs0 <= la_input[1];
	multiregimpl4_regs1 <= multiregimpl4_regs0;
	multiregimpl5_regs0 <= la_input[2];
	multiregimpl5_regs1 <= multiregimpl5_regs0;
	multiregimpl6_regs0 <= la_input[3];
	multiregimpl6_regs1 <= multiregimpl6_regs0;
	multiregimpl7_regs0 <= la_input[4];
	multiregimpl7_regs1 <= multiregimpl7_regs0;
	multiregimpl8_regs0 <= la_input[5];
	multiregimpl8_regs1 <= multiregimpl8_regs0;
	multiregimpl9_regs0 <= la_input[6];
	multiregimpl9_regs1 <= multiregimpl9_regs0;
	multiregimpl10_regs0 <= la_input[7];
	multiregimpl10_regs1 <= multiregimpl10_regs0;
	multiregimpl11_regs0 <= la_input[8];
	multiregimpl11_regs1 <= multiregimpl11_regs0;
	multiregimpl12_regs0 <= la_input[9];
	multiregimpl12_regs1 <= multiregimpl12_regs0;
	multiregimpl13_regs0 <= la_input[10];
	multiregimpl13_regs1 <= multiregimpl13_regs0;
	multiregimpl14_regs0 <= la_input[11];
	multiregimpl14_regs1 <= multiregimpl14_regs0;
	multiregimpl15_regs0 <= la_input[12];
	multiregimpl15_regs1 <= multiregimpl15_regs0;
	multiregimpl16_regs0 <= la_input[13];
	multiregimpl16_regs1 <= multiregimpl16_regs0;
	multiregimpl17_regs0 <= la_input[14];
	multiregimpl17_regs1 <= multiregimpl17_regs0;
	multiregimpl18_regs0 <= la_input[15];
	multiregimpl18_regs1 <= multiregimpl18_regs0;
	multiregimpl19_regs0 <= la_input[16];
	multiregimpl19_regs1 <= multiregimpl19_regs0;
	multiregimpl20_regs0 <= la_input[17];
	multiregimpl20_regs1 <= multiregimpl20_regs0;
	multiregimpl21_regs0 <= la_input[18];
	multiregimpl21_regs1 <= multiregimpl21_regs0;
	multiregimpl22_regs0 <= la_input[19];
	multiregimpl22_regs1 <= multiregimpl22_regs0;
	multiregimpl23_regs0 <= la_input[20];
	multiregimpl23_regs1 <= multiregimpl23_regs0;
	multiregimpl24_regs0 <= la_input[21];
	multiregimpl24_regs1 <= multiregimpl24_regs0;
	multiregimpl25_regs0 <= la_input[22];
	multiregimpl25_regs1 <= multiregimpl25_regs0;
	multiregimpl26_regs0 <= la_input[23];
	multiregimpl26_regs1 <= multiregimpl26_regs0;
	multiregimpl27_regs0 <= la_input[24];
	multiregimpl27_regs1 <= multiregimpl27_regs0;
	multiregimpl28_regs0 <= la_input[25];
	multiregimpl28_regs1 <= multiregimpl28_regs0;
	multiregimpl29_regs0 <= la_input[26];
	multiregimpl29_regs1 <= multiregimpl29_regs0;
	multiregimpl30_regs0 <= la_input[27];
	multiregimpl30_regs1 <= multiregimpl30_regs0;
	multiregimpl31_regs0 <= la_input[28];
	multiregimpl31_regs1 <= multiregimpl31_regs0;
	multiregimpl32_regs0 <= la_input[29];
	multiregimpl32_regs1 <= multiregimpl32_regs0;
	multiregimpl33_regs0 <= la_input[30];
	multiregimpl33_regs1 <= multiregimpl33_regs0;
	multiregimpl34_regs0 <= la_input[31];
	multiregimpl34_regs1 <= multiregimpl34_regs0;
	multiregimpl35_regs0 <= la_input[32];
	multiregimpl35_regs1 <= multiregimpl35_regs0;
	multiregimpl36_regs0 <= la_input[33];
	multiregimpl36_regs1 <= multiregimpl36_regs0;
	multiregimpl37_regs0 <= la_input[34];
	multiregimpl37_regs1 <= multiregimpl37_regs0;
	multiregimpl38_regs0 <= la_input[35];
	multiregimpl38_regs1 <= multiregimpl38_regs0;
	multiregimpl39_regs0 <= la_input[36];
	multiregimpl39_regs1 <= multiregimpl39_regs0;
	multiregimpl40_regs0 <= la_input[37];
	multiregimpl40_regs1 <= multiregimpl40_regs0;
	multiregimpl41_regs0 <= la_input[38];
	multiregimpl41_regs1 <= multiregimpl41_regs0;
	multiregimpl42_regs0 <= la_input[39];
	multiregimpl42_regs1 <= multiregimpl42_regs0;
	multiregimpl43_regs0 <= la_input[40];
	multiregimpl43_regs1 <= multiregimpl43_regs0;
	multiregimpl44_regs0 <= la_input[41];
	multiregimpl44_regs1 <= multiregimpl44_regs0;
	multiregimpl45_regs0 <= la_input[42];
	multiregimpl45_regs1 <= multiregimpl45_regs0;
	multiregimpl46_regs0 <= la_input[43];
	multiregimpl46_regs1 <= multiregimpl46_regs0;
	multiregimpl47_regs0 <= la_input[44];
	multiregimpl47_regs1 <= multiregimpl47_regs0;
	multiregimpl48_regs0 <= la_input[45];
	multiregimpl48_regs1 <= multiregimpl48_regs0;
	multiregimpl49_regs0 <= la_input[46];
	multiregimpl49_regs1 <= multiregimpl49_regs0;
	multiregimpl50_regs0 <= la_input[47];
	multiregimpl50_regs1 <= multiregimpl50_regs0;
	multiregimpl51_regs0 <= la_input[48];
	multiregimpl51_regs1 <= multiregimpl51_regs0;
	multiregimpl52_regs0 <= la_input[49];
	multiregimpl52_regs1 <= multiregimpl52_regs0;
	multiregimpl53_regs0 <= la_input[50];
	multiregimpl53_regs1 <= multiregimpl53_regs0;
	multiregimpl54_regs0 <= la_input[51];
	multiregimpl54_regs1 <= multiregimpl54_regs0;
	multiregimpl55_regs0 <= la_input[52];
	multiregimpl55_regs1 <= multiregimpl55_regs0;
	multiregimpl56_regs0 <= la_input[53];
	multiregimpl56_regs1 <= multiregimpl56_regs0;
	multiregimpl57_regs0 <= la_input[54];
	multiregimpl57_regs1 <= multiregimpl57_regs0;
	multiregimpl58_regs0 <= la_input[55];
	multiregimpl58_regs1 <= multiregimpl58_regs0;
	multiregimpl59_regs0 <= la_input[56];
	multiregimpl59_regs1 <= multiregimpl59_regs0;
	multiregimpl60_regs0 <= la_input[57];
	multiregimpl60_regs1 <= multiregimpl60_regs0;
	multiregimpl61_regs0 <= la_input[58];
	multiregimpl61_regs1 <= multiregimpl61_regs0;
	multiregimpl62_regs0 <= la_input[59];
	multiregimpl62_regs1 <= multiregimpl62_regs0;
	multiregimpl63_regs0 <= la_input[60];
	multiregimpl63_regs1 <= multiregimpl63_regs0;
	multiregimpl64_regs0 <= la_input[61];
	multiregimpl64_regs1 <= multiregimpl64_regs0;
	multiregimpl65_regs0 <= la_input[62];
	multiregimpl65_regs1 <= multiregimpl65_regs0;
	multiregimpl66_regs0 <= la_input[63];
	multiregimpl66_regs1 <= multiregimpl66_regs0;
	multiregimpl67_regs0 <= la_input[64];
	multiregimpl67_regs1 <= multiregimpl67_regs0;
	multiregimpl68_regs0 <= la_input[65];
	multiregimpl68_regs1 <= multiregimpl68_regs0;
	multiregimpl69_regs0 <= la_input[66];
	multiregimpl69_regs1 <= multiregimpl69_regs0;
	multiregimpl70_regs0 <= la_input[67];
	multiregimpl70_regs1 <= multiregimpl70_regs0;
	multiregimpl71_regs0 <= la_input[68];
	multiregimpl71_regs1 <= multiregimpl71_regs0;
	multiregimpl72_regs0 <= la_input[69];
	multiregimpl72_regs1 <= multiregimpl72_regs0;
	multiregimpl73_regs0 <= la_input[70];
	multiregimpl73_regs1 <= multiregimpl73_regs0;
	multiregimpl74_regs0 <= la_input[71];
	multiregimpl74_regs1 <= multiregimpl74_regs0;
	multiregimpl75_regs0 <= la_input[72];
	multiregimpl75_regs1 <= multiregimpl75_regs0;
	multiregimpl76_regs0 <= la_input[73];
	multiregimpl76_regs1 <= multiregimpl76_regs0;
	multiregimpl77_regs0 <= la_input[74];
	multiregimpl77_regs1 <= multiregimpl77_regs0;
	multiregimpl78_regs0 <= la_input[75];
	multiregimpl78_regs1 <= multiregimpl78_regs0;
	multiregimpl79_regs0 <= la_input[76];
	multiregimpl79_regs1 <= multiregimpl79_regs0;
	multiregimpl80_regs0 <= la_input[77];
	multiregimpl80_regs1 <= multiregimpl80_regs0;
	multiregimpl81_regs0 <= la_input[78];
	multiregimpl81_regs1 <= multiregimpl81_regs0;
	multiregimpl82_regs0 <= la_input[79];
	multiregimpl82_regs1 <= multiregimpl82_regs0;
	multiregimpl83_regs0 <= la_input[80];
	multiregimpl83_regs1 <= multiregimpl83_regs0;
	multiregimpl84_regs0 <= la_input[81];
	multiregimpl84_regs1 <= multiregimpl84_regs0;
	multiregimpl85_regs0 <= la_input[82];
	multiregimpl85_regs1 <= multiregimpl85_regs0;
	multiregimpl86_regs0 <= la_input[83];
	multiregimpl86_regs1 <= multiregimpl86_regs0;
	multiregimpl87_regs0 <= la_input[84];
	multiregimpl87_regs1 <= multiregimpl87_regs0;
	multiregimpl88_regs0 <= la_input[85];
	multiregimpl88_regs1 <= multiregimpl88_regs0;
	multiregimpl89_regs0 <= la_input[86];
	multiregimpl89_regs1 <= multiregimpl89_regs0;
	multiregimpl90_regs0 <= la_input[87];
	multiregimpl90_regs1 <= multiregimpl90_regs0;
	multiregimpl91_regs0 <= la_input[88];
	multiregimpl91_regs1 <= multiregimpl91_regs0;
	multiregimpl92_regs0 <= la_input[89];
	multiregimpl92_regs1 <= multiregimpl92_regs0;
	multiregimpl93_regs0 <= la_input[90];
	multiregimpl93_regs1 <= multiregimpl93_regs0;
	multiregimpl94_regs0 <= la_input[91];
	multiregimpl94_regs1 <= multiregimpl94_regs0;
	multiregimpl95_regs0 <= la_input[92];
	multiregimpl95_regs1 <= multiregimpl95_regs0;
	multiregimpl96_regs0 <= la_input[93];
	multiregimpl96_regs1 <= multiregimpl96_regs0;
	multiregimpl97_regs0 <= la_input[94];
	multiregimpl97_regs1 <= multiregimpl97_regs0;
	multiregimpl98_regs0 <= la_input[95];
	multiregimpl98_regs1 <= multiregimpl98_regs0;
	multiregimpl99_regs0 <= la_input[96];
	multiregimpl99_regs1 <= multiregimpl99_regs0;
	multiregimpl100_regs0 <= la_input[97];
	multiregimpl100_regs1 <= multiregimpl100_regs0;
	multiregimpl101_regs0 <= la_input[98];
	multiregimpl101_regs1 <= multiregimpl101_regs0;
	multiregimpl102_regs0 <= la_input[99];
	multiregimpl102_regs1 <= multiregimpl102_regs0;
	multiregimpl103_regs0 <= la_input[100];
	multiregimpl103_regs1 <= multiregimpl103_regs0;
	multiregimpl104_regs0 <= la_input[101];
	multiregimpl104_regs1 <= multiregimpl104_regs0;
	multiregimpl105_regs0 <= la_input[102];
	multiregimpl105_regs1 <= multiregimpl105_regs0;
	multiregimpl106_regs0 <= la_input[103];
	multiregimpl106_regs1 <= multiregimpl106_regs0;
	multiregimpl107_regs0 <= la_input[104];
	multiregimpl107_regs1 <= multiregimpl107_regs0;
	multiregimpl108_regs0 <= la_input[105];
	multiregimpl108_regs1 <= multiregimpl108_regs0;
	multiregimpl109_regs0 <= la_input[106];
	multiregimpl109_regs1 <= multiregimpl109_regs0;
	multiregimpl110_regs0 <= la_input[107];
	multiregimpl110_regs1 <= multiregimpl110_regs0;
	multiregimpl111_regs0 <= la_input[108];
	multiregimpl111_regs1 <= multiregimpl111_regs0;
	multiregimpl112_regs0 <= la_input[109];
	multiregimpl112_regs1 <= multiregimpl112_regs0;
	multiregimpl113_regs0 <= la_input[110];
	multiregimpl113_regs1 <= multiregimpl113_regs0;
	multiregimpl114_regs0 <= la_input[111];
	multiregimpl114_regs1 <= multiregimpl114_regs0;
	multiregimpl115_regs0 <= la_input[112];
	multiregimpl115_regs1 <= multiregimpl115_regs0;
	multiregimpl116_regs0 <= la_input[113];
	multiregimpl116_regs1 <= multiregimpl116_regs0;
	multiregimpl117_regs0 <= la_input[114];
	multiregimpl117_regs1 <= multiregimpl117_regs0;
	multiregimpl118_regs0 <= la_input[115];
	multiregimpl118_regs1 <= multiregimpl118_regs0;
	multiregimpl119_regs0 <= la_input[116];
	multiregimpl119_regs1 <= multiregimpl119_regs0;
	multiregimpl120_regs0 <= la_input[117];
	multiregimpl120_regs1 <= multiregimpl120_regs0;
	multiregimpl121_regs0 <= la_input[118];
	multiregimpl121_regs1 <= multiregimpl121_regs0;
	multiregimpl122_regs0 <= la_input[119];
	multiregimpl122_regs1 <= multiregimpl122_regs0;
	multiregimpl123_regs0 <= la_input[120];
	multiregimpl123_regs1 <= multiregimpl123_regs0;
	multiregimpl124_regs0 <= la_input[121];
	multiregimpl124_regs1 <= multiregimpl124_regs0;
	multiregimpl125_regs0 <= la_input[122];
	multiregimpl125_regs1 <= multiregimpl125_regs0;
	multiregimpl126_regs0 <= la_input[123];
	multiregimpl126_regs1 <= multiregimpl126_regs0;
	multiregimpl127_regs0 <= la_input[124];
	multiregimpl127_regs1 <= multiregimpl127_regs0;
	multiregimpl128_regs0 <= la_input[125];
	multiregimpl128_regs1 <= multiregimpl128_regs0;
	multiregimpl129_regs0 <= la_input[126];
	multiregimpl129_regs1 <= multiregimpl129_regs0;
	multiregimpl130_regs0 <= la_input[127];
	multiregimpl130_regs1 <= multiregimpl130_regs0;
	multiregimpl131_regs0 <= user_irq[0];
	multiregimpl131_regs1 <= multiregimpl131_regs0;
	multiregimpl132_regs0 <= user_irq[1];
	multiregimpl132_regs1 <= multiregimpl132_regs0;
	multiregimpl133_regs0 <= user_irq[2];
	multiregimpl133_regs1 <= multiregimpl133_regs0;
	multiregimpl134_regs0 <= user_irq[3];
	multiregimpl134_regs1 <= multiregimpl134_regs0;
	multiregimpl135_regs0 <= user_irq[4];
	multiregimpl135_regs1 <= multiregimpl135_regs0;
	multiregimpl136_regs0 <= user_irq[5];
	multiregimpl136_regs1 <= multiregimpl136_regs0;
end

RAM256 RAM256(
	.A0(dff_bus_adr[7:0]),
	.CLK(sys_clk),
	.Di0(dff_di),
	.EN0(dff_en),
	.WE0(dff_we),
	.Do0(dff_do)
);

RAM128 RAM128(
	.A0(dff2_bus_adr[6:0]),
	.CLK(sys_clk),
	.Di0(dff2_di),
	.EN0(dff2_en),
	.WE0(dff2_we),
	.Do0(dff2_do)
);

reg [9:0] storage[0:15];
reg [9:0] memdat;
reg [9:0] memdat_1;
always @(posedge sys_clk) begin
	if (uart_tx_fifo_wrport_we)
		storage[uart_tx_fifo_wrport_adr] <= uart_tx_fifo_wrport_dat_w;
	memdat <= storage[uart_tx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (uart_tx_fifo_rdport_re)
		memdat_1 <= storage[uart_tx_fifo_rdport_adr];
end

assign uart_tx_fifo_wrport_dat_r = memdat;
assign uart_tx_fifo_rdport_dat_r = memdat_1;

reg [9:0] storage_1[0:15];
reg [9:0] memdat_2;
reg [9:0] memdat_3;
always @(posedge sys_clk) begin
	if (uart_rx_fifo_wrport_we)
		storage_1[uart_rx_fifo_wrport_adr] <= uart_rx_fifo_wrport_dat_w;
	memdat_2 <= storage_1[uart_rx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (uart_rx_fifo_rdport_re)
		memdat_3 <= storage_1[uart_rx_fifo_rdport_adr];
end

assign uart_rx_fifo_wrport_dat_r = memdat_2;
assign uart_rx_fifo_rdport_dat_r = memdat_3;

VexRiscv VexRiscv(

    .vccd1(VPWR),
    .vssd1(VGND),

	.clk(sys_clk),
	.dBusWishbone_ACK(mgmtsoc_dbus_dbus_ack),
	.dBusWishbone_DAT_MISO(mgmtsoc_dbus_dbus_dat_r),
	.dBusWishbone_ERR((mgmtsoc_dbus_dbus_err | mgmtsoc_vexriscv_dbus_err)),
	.debugReset(sys_rst),
	.debug_bus_cmd_payload_address(mgmtsoc_vexriscv_i_cmd_payload_address),
	.debug_bus_cmd_payload_data(mgmtsoc_vexriscv_i_cmd_payload_data),
	.debug_bus_cmd_payload_wr(mgmtsoc_vexriscv_i_cmd_payload_wr),
	.debug_bus_cmd_valid(mgmtsoc_vexriscv_i_cmd_valid),
	.externalInterruptArray(mgmtsoc_interrupt),
	.externalResetVector(mgmtsoc_vexriscv),
	.iBusWishbone_ACK(mgmtsoc_ibus_ibus_ack),
	.iBusWishbone_DAT_MISO(mgmtsoc_ibus_ibus_dat_r),
	.iBusWishbone_ERR((mgmtsoc_ibus_ibus_err | mgmtsoc_vexriscv_ibus_err)),
	.reset(((sys_rst | mgmtsoc_reset) | mgmtsoc_vexriscv_debug_reset)),
	.softwareInterrupt(1'd0),
	.timerInterrupt(1'd0),
	.dBusWishbone_ADR(mgmtsoc_dbus_dbus_adr),
	.dBusWishbone_BTE(mgmtsoc_dbus_dbus_bte),
	.dBusWishbone_CTI(mgmtsoc_dbus_dbus_cti),
	.dBusWishbone_CYC(mgmtsoc_dbus_dbus_cyc),
	.dBusWishbone_DAT_MOSI(mgmtsoc_dbus_dbus_dat_w),
	.dBusWishbone_SEL(mgmtsoc_dbus_dbus_sel),
	.dBusWishbone_STB(mgmtsoc_dbus_dbus_stb),
	.dBusWishbone_WE(mgmtsoc_dbus_dbus_we),
	.debug_bus_cmd_ready(mgmtsoc_vexriscv_o_cmd_ready),
	.debug_bus_rsp_data(mgmtsoc_vexriscv_o_rsp_data),
	.debug_resetOut(mgmtsoc_vexriscv_o_resetOut),
	.iBusWishbone_ADR(mgmtsoc_ibus_ibus_adr),
	.iBusWishbone_BTE(mgmtsoc_ibus_ibus_bte),
	.iBusWishbone_CTI(mgmtsoc_ibus_ibus_cti),
	.iBusWishbone_CYC(mgmtsoc_ibus_ibus_cyc),
	.iBusWishbone_DAT_MOSI(mgmtsoc_ibus_ibus_dat_w),
	.iBusWishbone_SEL(mgmtsoc_ibus_ibus_sel),
	.iBusWishbone_STB(mgmtsoc_ibus_ibus_stb),
	.iBusWishbone_WE(mgmtsoc_ibus_ibus_we)
);

endmodule
/*
 *  SPDX-FileCopyrightText: 2015 Clifford Wolf
 *  PicoSoC - A simple example SoC using PicoRV32
 *
 *  Copyright (C) 2017  Clifford Wolf <clifford@clifford.at>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 *  Revision 1,  July 2019:  Added signals to drive flash_clk and flash_csb
 *  output enable (inverted), tied to reset so that the flash is completely
 *  isolated from the processor when the processor is in reset.
 *
 *  Also: Made ram_wenb a 4-bit bus so that the memory access can be made
 *  byte-wide for byte-wide instructions.
 *
 *  SPDX-License-Identifier: ISC
 */


`default_nettype none




/* Wrapper module around management SoC core for pin compatibility  */
/* with the Caravel harness chip. */    

module mgmt_core_wrapper (

    inout VPWR,     /* 1.8V domain */
    inout VGND,

    // Clock and reset
    input core_clk,
    input core_rstn,

    // GPIO (one pin)
    output gpio_out_pad,    // Connect to out on gpio pad
    input  gpio_in_pad,     // Connect to in on gpio pad
    output gpio_mode0_pad,  // Connect to dm[0] on gpio pad
    output gpio_mode1_pad,  // Connect to dm[2] on gpio pad
    output gpio_outenb_pad, // Connect to oe_n on gpio pad
    output gpio_inenb_pad,  // Connect to inp_dis on gpio pad

    // Logic analyzer signals
    input  [127:0] la_input,            // From user project to CPU
    output [127:0] la_output,           // From CPU to user project
    output [127:0] la_oenb,             // Logic analyzer output enable
    output [127:0] la_iena,             // Logic analyzer input enable

    // Flash memory control (SPI master)
    output flash_csb,
    output flash_clk,

    output flash_io0_oeb,
    output flash_io1_oeb,
    output flash_io2_oeb,
    output flash_io3_oeb,

    output flash_io0_do,
    output flash_io1_do,
    output flash_io2_do,
    output flash_io3_do,

    input  flash_io0_di,
    input  flash_io1_di,
    input  flash_io2_di,
    input  flash_io3_di,

    // Exported Wishboned bus
    output    mprj_wb_iena, // Enable for the user wishbone return signals
    output    mprj_cyc_o,
    output    mprj_stb_o,
    output    mprj_we_o,
    output [3:0]  mprj_sel_o,
    output [31:0] mprj_adr_o,
    output [31:0] mprj_dat_o,
    input     mprj_ack_i,
    input  [31:0] mprj_dat_i,

    output    hk_cyc_o,
    output    hk_stb_o,
    input  [31:0] hk_dat_i,
    input     hk_ack_i,

    // IRQ
    input  [5:0] irq,       // IRQ from SPI and user project
    output [2:0] user_irq_ena,  // Enables for user project IRQ

    // Module status
    output qspi_enabled,
    output uart_enabled,
    output spi_enabled,
    output debug_mode,

    // Module I/O
    output ser_tx,
    input  ser_rx,
    output spi_csb,
    output spi_sck,
    output spi_sdo,
    output spi_sdoenb,
    input  spi_sdi,
    input  debug_in,
    output debug_out,
    output debug_oeb,

    // Trap state from CPU
    output trap
);


// Signals below are sram_ro ports that left no_connect
// as they are tied down inside mgmt_core

    /* Implement the PicoSoC core */

    mgmt_core core (
    
        .VPWR(VPWR),        /* 1.8V domain */
        .VGND(VGND),
    
        .core_clk(core_clk),
        .core_rstn(core_rstn),

        // Trap state from CPU
        .trap(trap),

        // GPIO (one pin)
        .gpio_out_pad(gpio_out_pad),        // Connect to out on gpio pad
        .gpio_in_pad(gpio_in_pad),      // Connect to in on gpio pad
        .gpio_mode0_pad(gpio_mode0_pad),    // Connect to dm[0] on gpio pad
        .gpio_mode1_pad(gpio_mode1_pad),    // Connect to dm[2] on gpio pad
        .gpio_outenb_pad(gpio_outenb_pad),  // Connect to oe_n on gpio pad
        .gpio_inenb_pad(gpio_inenb_pad),    // Connect to inp_dis on gpio pad

        .la_input(la_input),            // From user project to CPU
        .la_output(la_output),          // From CPU to user project
        .la_oenb(la_oenb),          // Logic analyzer output enable
        .la_iena(la_iena),          // Logic analyzer input enable

        // IRQ
        .user_irq(irq),     // IRQ from SPI and user project
        .user_irq_ena(user_irq_ena),

        // Flash memory control (SPI master)
        .flash_cs_n(flash_csb),
        .flash_clk(flash_clk),

        .flash_io0_oeb(flash_io0_oeb),
        .flash_io1_oeb(flash_io1_oeb),
        .flash_io2_oeb(flash_io2_oeb),
        .flash_io3_oeb(flash_io3_oeb),

        .flash_io0_do(flash_io0_do),
        .flash_io1_do(flash_io1_do),
        .flash_io2_do(flash_io2_do),
        .flash_io3_do(flash_io3_do),

        .flash_io0_di(flash_io0_di),
        .flash_io1_di(flash_io1_di),
        .flash_io2_di(flash_io2_di),
        .flash_io3_di(flash_io3_di),

        // Exported wishbone bus (User project)
        .mprj_wb_iena(mprj_wb_iena),
        .mprj_ack_i(mprj_ack_i),
        .mprj_dat_i(mprj_dat_i),
        .mprj_cyc_o(mprj_cyc_o),
        .mprj_stb_o(mprj_stb_o),
        .mprj_we_o(mprj_we_o),
        .mprj_sel_o(mprj_sel_o),
        .mprj_adr_o(mprj_adr_o),
        .mprj_dat_o(mprj_dat_o),

        .hk_cyc_o(hk_cyc_o),
        .hk_stb_o(hk_stb_o),
        .hk_dat_i(hk_dat_i),
        .hk_ack_i(hk_ack_i),

        // Module status
        .qspi_enabled(qspi_enabled),
        .uart_enabled(uart_enabled),
        .spi_enabled(spi_enabled),
        .debug_mode(debug_mode),

        // Module I/O
//      .ser_tx(ser_tx),
//      .ser_rx(ser_rx),
        .serial_tx(ser_tx),
        .serial_rx(ser_rx),
        .spi_cs_n(spi_csb),
        .spi_clk(spi_sck),
        .spi_miso(spi_sdi),
        .spi_sdoenb(spi_sdoenb),
        .spi_mosi(spi_sdo),
        .debug_in(debug_in),
        .debug_out(debug_out),
        .debug_oeb(debug_oeb)

    );


endmodule
`default_nettype wire


// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : VexRiscv
// Git hash  : c4eca1837ebca20b637a0a61e3a93d9446488459










































module VexRiscv (

    inout vccd1,	    /* 1.8V domain */
    inout vssd1,

  input      [31:0]   externalResetVector,
  input               timerInterrupt,
  input               softwareInterrupt,
  input      [31:0]   externalInterruptArray,
  input               debug_bus_cmd_valid,
  output reg          debug_bus_cmd_ready,
  input               debug_bus_cmd_payload_wr,
  input      [7:0]    debug_bus_cmd_payload_address,
  input      [31:0]   debug_bus_cmd_payload_data,
  output reg [31:0]   debug_bus_rsp_data,
  output              debug_resetOut,
  output reg          iBusWishbone_CYC,
  output reg          iBusWishbone_STB,
  input               iBusWishbone_ACK,
  output              iBusWishbone_WE,
  output     [29:0]   iBusWishbone_ADR,
  input      [31:0]   iBusWishbone_DAT_MISO,
  output     [31:0]   iBusWishbone_DAT_MOSI,
  output     [3:0]    iBusWishbone_SEL,
  input               iBusWishbone_ERR,
  output     [2:0]    iBusWishbone_CTI,
  output     [1:0]    iBusWishbone_BTE,
  output              dBusWishbone_CYC,
  output              dBusWishbone_STB,
  input               dBusWishbone_ACK,
  output              dBusWishbone_WE,
  output     [29:0]   dBusWishbone_ADR,
  input      [31:0]   dBusWishbone_DAT_MISO,
  output     [31:0]   dBusWishbone_DAT_MOSI,
  output reg [3:0]    dBusWishbone_SEL,
  input               dBusWishbone_ERR,
  output     [2:0]    dBusWishbone_CTI,
  output     [1:0]    dBusWishbone_BTE,
  input               clk,
  input               reset,
  input               debugReset
);
  wire                IBusCachedPlugin_cache_io_flush;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isRemoved;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isUser;
  reg                 IBusCachedPlugin_cache_io_cpu_fill_valid;
  reg        [31:0]   _zz_RegFilePlugin_regFile_port0;
  reg        [31:0]   _zz_RegFilePlugin_regFile_port1;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_haltIt;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_data;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress;
  wire                IBusCachedPlugin_cache_io_cpu_decode_error;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuException;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_data;
  wire                IBusCachedPlugin_cache_io_cpu_decode_cacheMiss;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_physicalAddress;
  wire                IBusCachedPlugin_cache_io_mem_cmd_valid;
  wire       [31:0]   IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  wire       [2:0]    IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_1;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_2;
  wire                _zz_decode_LEGAL_INSTRUCTION_3;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_4;
  wire       [12:0]   _zz_decode_LEGAL_INSTRUCTION_5;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_6;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_7;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_8;
  wire                _zz_decode_LEGAL_INSTRUCTION_9;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_10;
  wire       [6:0]    _zz_decode_LEGAL_INSTRUCTION_11;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_12;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_13;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_14;
  wire                _zz_decode_LEGAL_INSTRUCTION_15;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_16;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_17;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_1;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_2;
  wire       [31:0]   _zz_IBusCachedPlugin_fetchPc_pc;
  wire       [2:0]    _zz_IBusCachedPlugin_fetchPc_pc_1;
  wire       [2:0]    _zz_DBusSimplePlugin_memoryExceptionPort_payload_code;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_1;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_2;
  wire                _zz__zz_decode_ENV_CTRL_2_3;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_4;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_5;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_6;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_7;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_8;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_9;
  wire                _zz__zz_decode_ENV_CTRL_2_10;
  wire                _zz__zz_decode_ENV_CTRL_2_11;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_12;
  wire                _zz__zz_decode_ENV_CTRL_2_13;
  wire       [21:0]   _zz__zz_decode_ENV_CTRL_2_14;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_15;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_16;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_17;
  wire                _zz__zz_decode_ENV_CTRL_2_18;
  wire                _zz__zz_decode_ENV_CTRL_2_19;
  wire                _zz__zz_decode_ENV_CTRL_2_20;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_21;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_22;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_23;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_24;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_25;
  wire       [18:0]   _zz__zz_decode_ENV_CTRL_2_26;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_27;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_28;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_29;
  wire                _zz__zz_decode_ENV_CTRL_2_30;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_31;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_32;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_33;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_34;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_35;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_36;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_37;
  wire       [15:0]   _zz__zz_decode_ENV_CTRL_2_38;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_39;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_40;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_41;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_42;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_43;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_44;
  wire                _zz__zz_decode_ENV_CTRL_2_45;
  wire                _zz__zz_decode_ENV_CTRL_2_46;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_47;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_48;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_49;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_50;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_51;
  wire                _zz__zz_decode_ENV_CTRL_2_52;
  wire       [12:0]   _zz__zz_decode_ENV_CTRL_2_53;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_54;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_55;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_56;
  wire                _zz__zz_decode_ENV_CTRL_2_57;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_58;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_59;
  wire       [4:0]    _zz__zz_decode_ENV_CTRL_2_60;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_61;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_62;
  wire                _zz__zz_decode_ENV_CTRL_2_63;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_64;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_65;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_66;
  wire                _zz__zz_decode_ENV_CTRL_2_67;
  wire                _zz__zz_decode_ENV_CTRL_2_68;
  wire       [9:0]    _zz__zz_decode_ENV_CTRL_2_69;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_70;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_71;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_72;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_73;
  wire                _zz__zz_decode_ENV_CTRL_2_74;
  wire                _zz__zz_decode_ENV_CTRL_2_75;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_76;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_77;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_78;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_79;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_80;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_81;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_82;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_83;
  wire       [6:0]    _zz__zz_decode_ENV_CTRL_2_84;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_85;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_86;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_87;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_88;
  wire                _zz__zz_decode_ENV_CTRL_2_89;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_90;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_91;
  wire       [2:0]    _zz__zz_decode_ENV_CTRL_2_92;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_93;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_94;
  wire                _zz__zz_decode_ENV_CTRL_2_95;
  wire                _zz__zz_decode_ENV_CTRL_2_96;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_97;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_98;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_99;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_100;
  wire       [3:0]    _zz__zz_decode_ENV_CTRL_2_101;
  wire                _zz__zz_decode_ENV_CTRL_2_102;
  wire                _zz__zz_decode_ENV_CTRL_2_103;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_104;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_105;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_106;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_107;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_108;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_109;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_110;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_111;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_112;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_113;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_114;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_115;
  wire       [1:0]    _zz__zz_decode_ENV_CTRL_2_116;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_117;
  wire       [31:0]   _zz__zz_decode_ENV_CTRL_2_118;
  wire       [0:0]    _zz__zz_decode_ENV_CTRL_2_119;
  wire                _zz_RegFilePlugin_regFile_port;
  wire                _zz_decode_RegFilePlugin_rs1Data;
  wire                _zz_RegFilePlugin_regFile_port_1;
  wire                _zz_decode_RegFilePlugin_rs2Data;
  wire       [0:0]    _zz__zz_execute_REGFILE_WRITE_DATA;
  wire       [2:0]    _zz__zz_execute_SRC1;
  wire       [4:0]    _zz__zz_execute_SRC1_1;
  wire       [11:0]   _zz__zz_execute_SRC2_3;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_1;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_2;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_3;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_4;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_5;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_6;
  wire       [31:0]   _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1;
  wire       [32:0]   _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1_1;
  wire       [19:0]   _zz__zz_execute_BranchPlugin_branch_src2;
  wire       [11:0]   _zz__zz_execute_BranchPlugin_branch_src2_4;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3_1;
  wire                _zz_when;
  wire                _zz_when_1;
  wire       [26:0]   _zz_iBusWishbone_ADR_1;
  wire       [31:0]   memory_MEMORY_READ_DATA;
  wire       [31:0]   execute_BRANCH_CALC;
  wire                execute_BRANCH_DO;
  wire       [31:0]   writeBack_REGFILE_WRITE_DATA;
  wire       [31:0]   execute_REGFILE_WRITE_DATA;
  wire       [1:0]    memory_MEMORY_ADDRESS_LOW;
  wire       [1:0]    execute_MEMORY_ADDRESS_LOW;
  wire                decode_DO_EBREAK;
  wire                decode_CSR_READ_OPCODE;
  wire                decode_CSR_WRITE_OPCODE;
  wire                decode_SRC2_FORCE_ZERO;
  wire       [31:0]   decode_RS2;
  wire       [31:0]   decode_RS1;
  wire       [1:0] _zz_memory_to_writeBack_ENV_CTRL;
  wire       [1:0] _zz_memory_to_writeBack_ENV_CTRL_1;
  wire       [1:0] _zz_execute_to_memory_ENV_CTRL;
  wire       [1:0] _zz_execute_to_memory_ENV_CTRL_1;
  wire       [1:0] decode_ENV_CTRL;
  wire       [1:0] _zz_decode_ENV_CTRL;
  wire       [1:0] _zz_decode_to_execute_ENV_CTRL;
  wire       [1:0] _zz_decode_to_execute_ENV_CTRL_1;
  wire                decode_IS_CSR;
  wire       [1:0] decode_BRANCH_CTRL;
  wire       [1:0] _zz_decode_BRANCH_CTRL;
  wire       [1:0] _zz_decode_to_execute_BRANCH_CTRL;
  wire       [1:0] _zz_decode_to_execute_BRANCH_CTRL_1;
  wire       [1:0] decode_SHIFT_CTRL;
  wire       [1:0] _zz_decode_SHIFT_CTRL;
  wire       [1:0] _zz_decode_to_execute_SHIFT_CTRL;
  wire       [1:0] _zz_decode_to_execute_SHIFT_CTRL_1;
  wire       [1:0] decode_ALU_BITWISE_CTRL;
  wire       [1:0] _zz_decode_ALU_BITWISE_CTRL;
  wire       [1:0] _zz_decode_to_execute_ALU_BITWISE_CTRL;
  wire       [1:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  wire                decode_SRC_LESS_UNSIGNED;
  wire                decode_MEMORY_STORE;
  wire                execute_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_EXECUTE_STAGE;
  wire       [1:0] decode_SRC2_CTRL;
  wire       [1:0] _zz_decode_SRC2_CTRL;
  wire       [1:0] _zz_decode_to_execute_SRC2_CTRL;
  wire       [1:0] _zz_decode_to_execute_SRC2_CTRL_1;
  wire       [1:0] decode_ALU_CTRL;
  wire       [1:0] _zz_decode_ALU_CTRL;
  wire       [1:0] _zz_decode_to_execute_ALU_CTRL;
  wire       [1:0] _zz_decode_to_execute_ALU_CTRL_1;
  wire                decode_MEMORY_ENABLE;
  wire       [1:0] decode_SRC1_CTRL;
  wire       [1:0] _zz_decode_SRC1_CTRL;
  wire       [1:0] _zz_decode_to_execute_SRC1_CTRL;
  wire       [1:0] _zz_decode_to_execute_SRC1_CTRL_1;
  wire       [31:0]   writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   memory_FORMAL_PC_NEXT;
  wire       [31:0]   execute_FORMAL_PC_NEXT;
  wire       [31:0]   decode_FORMAL_PC_NEXT;
  wire       [31:0]   memory_PC;
  wire                execute_DO_EBREAK;
  wire                decode_IS_EBREAK;
  wire                execute_CSR_READ_OPCODE;
  wire                execute_CSR_WRITE_OPCODE;
  wire                execute_IS_CSR;
  wire       [1:0] memory_ENV_CTRL;
  wire       [1:0] _zz_memory_ENV_CTRL;
  wire       [1:0] execute_ENV_CTRL;
  wire       [1:0] _zz_execute_ENV_CTRL;
  wire       [1:0] writeBack_ENV_CTRL;
  wire       [1:0] _zz_writeBack_ENV_CTRL;
  wire       [31:0]   memory_BRANCH_CALC;
  wire                memory_BRANCH_DO;
  wire       [31:0]   execute_PC;
  wire       [31:0]   execute_RS1;
  wire       [1:0] execute_BRANCH_CTRL;
  wire       [1:0] _zz_execute_BRANCH_CTRL;
  wire                decode_RS2_USE;
  wire                decode_RS1_USE;
  wire                execute_REGFILE_WRITE_VALID;
  wire                execute_BYPASSABLE_EXECUTE_STAGE;
  wire                memory_REGFILE_WRITE_VALID;
  wire       [31:0]   memory_INSTRUCTION;
  wire                memory_BYPASSABLE_MEMORY_STAGE;
  wire                writeBack_REGFILE_WRITE_VALID;
  reg        [31:0]   _zz_execute_to_memory_REGFILE_WRITE_DATA;
  wire       [1:0] execute_SHIFT_CTRL;
  wire       [1:0] _zz_execute_SHIFT_CTRL;
  wire                execute_SRC_LESS_UNSIGNED;
  wire                execute_SRC2_FORCE_ZERO;
  wire                execute_SRC_USE_SUB_LESS;
  wire       [31:0]   _zz_execute_SRC2;
  wire       [1:0] execute_SRC2_CTRL;
  wire       [1:0] _zz_execute_SRC2_CTRL;
  wire       [1:0] execute_SRC1_CTRL;
  wire       [1:0] _zz_execute_SRC1_CTRL;
  wire                decode_SRC_USE_SUB_LESS;
  wire                decode_SRC_ADD_ZERO;
  wire       [31:0]   execute_SRC_ADD_SUB;
  wire                execute_SRC_LESS;
  wire       [1:0] execute_ALU_CTRL;
  wire       [1:0] _zz_execute_ALU_CTRL;
  wire       [31:0]   execute_SRC2;
  wire       [31:0]   execute_SRC1;
  wire       [1:0] execute_ALU_BITWISE_CTRL;
  wire       [1:0] _zz_execute_ALU_BITWISE_CTRL;
  wire       [31:0]   _zz_lastStageRegFileWrite_payload_address;
  wire                _zz_lastStageRegFileWrite_valid;
  reg                 _zz_1;
  wire       [31:0]   decode_INSTRUCTION_ANTICIPATED;
  reg                 decode_REGFILE_WRITE_VALID;
  wire                decode_LEGAL_INSTRUCTION;
  wire       [1:0] _zz_decode_ENV_CTRL_1;
  wire       [1:0] _zz_decode_BRANCH_CTRL_1;
  wire       [1:0] _zz_decode_SHIFT_CTRL_1;
  wire       [1:0] _zz_decode_ALU_BITWISE_CTRL_1;
  wire       [1:0] _zz_decode_SRC2_CTRL_1;
  wire       [1:0] _zz_decode_ALU_CTRL_1;
  wire       [1:0] _zz_decode_SRC1_CTRL_1;
  wire                writeBack_MEMORY_STORE;
  reg        [31:0]   _zz_lastStageRegFileWrite_payload_data;
  wire                writeBack_MEMORY_ENABLE;
  wire       [1:0]    writeBack_MEMORY_ADDRESS_LOW;
  wire       [31:0]   writeBack_MEMORY_READ_DATA;
  wire                memory_ALIGNEMENT_FAULT;
  wire       [31:0]   memory_REGFILE_WRITE_DATA;
  wire                memory_MEMORY_STORE;
  wire                memory_MEMORY_ENABLE;
  wire       [31:0]   execute_SRC_ADD;
  wire       [31:0]   execute_RS2;
  wire       [31:0]   execute_INSTRUCTION;
  wire                execute_MEMORY_STORE;
  wire                execute_MEMORY_ENABLE;
  wire                execute_ALIGNEMENT_FAULT;
  wire                decode_FLUSH_ALL;
  reg                 IBusCachedPlugin_rsp_issueDetected_4;
  reg                 IBusCachedPlugin_rsp_issueDetected_3;
  reg                 IBusCachedPlugin_rsp_issueDetected_2;
  reg                 IBusCachedPlugin_rsp_issueDetected_1;
  wire       [31:0]   decode_INSTRUCTION;
  reg        [31:0]   _zz_memory_to_writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   decode_PC;
  wire       [31:0]   writeBack_PC;
  wire       [31:0]   writeBack_INSTRUCTION;
  reg                 decode_arbitration_haltItself;
  reg                 decode_arbitration_haltByOther;
  reg                 decode_arbitration_removeIt;
  wire                decode_arbitration_flushIt;
  reg                 decode_arbitration_flushNext;
  reg                 decode_arbitration_isValid;
  wire                decode_arbitration_isStuck;
  wire                decode_arbitration_isStuckByOthers;
  wire                decode_arbitration_isFlushed;
  wire                decode_arbitration_isMoving;
  wire                decode_arbitration_isFiring;
  reg                 execute_arbitration_haltItself;
  reg                 execute_arbitration_haltByOther;
  reg                 execute_arbitration_removeIt;
  reg                 execute_arbitration_flushIt;
  reg                 execute_arbitration_flushNext;
  reg                 execute_arbitration_isValid;
  wire                execute_arbitration_isStuck;
  wire                execute_arbitration_isStuckByOthers;
  wire                execute_arbitration_isFlushed;
  wire                execute_arbitration_isMoving;
  wire                execute_arbitration_isFiring;
  reg                 memory_arbitration_haltItself;
  wire                memory_arbitration_haltByOther;
  reg                 memory_arbitration_removeIt;
  wire                memory_arbitration_flushIt;
  reg                 memory_arbitration_flushNext;
  reg                 memory_arbitration_isValid;
  wire                memory_arbitration_isStuck;
  wire                memory_arbitration_isStuckByOthers;
  wire                memory_arbitration_isFlushed;
  wire                memory_arbitration_isMoving;
  wire                memory_arbitration_isFiring;
  wire                writeBack_arbitration_haltItself;
  wire                writeBack_arbitration_haltByOther;
  reg                 writeBack_arbitration_removeIt;
  wire                writeBack_arbitration_flushIt;
  reg                 writeBack_arbitration_flushNext;
  reg                 writeBack_arbitration_isValid;
  wire                writeBack_arbitration_isStuck;
  wire                writeBack_arbitration_isStuckByOthers;
  wire                writeBack_arbitration_isFlushed;
  wire                writeBack_arbitration_isMoving;
  wire                writeBack_arbitration_isFiring;
  wire       [31:0]   lastStageInstruction /* verilator public */ ;
  wire       [31:0]   lastStagePc /* verilator public */ ;
  wire                lastStageIsValid /* verilator public */ ;
  wire                lastStageIsFiring /* verilator public */ ;
  reg                 IBusCachedPlugin_fetcherHalt;
  reg                 IBusCachedPlugin_incomingInstruction;
  wire                IBusCachedPlugin_pcValids_0;
  wire                IBusCachedPlugin_pcValids_1;
  wire                IBusCachedPlugin_pcValids_2;
  wire                IBusCachedPlugin_pcValids_3;
  reg                 IBusCachedPlugin_decodeExceptionPort_valid;
  reg        [3:0]    IBusCachedPlugin_decodeExceptionPort_payload_code;
  wire       [31:0]   IBusCachedPlugin_decodeExceptionPort_payload_badAddr;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isValid;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isStuck;
  wire       [31:0]   IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  wire                IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation;
  wire       [31:0]   IBusCachedPlugin_mmuBus_rsp_physicalAddress;
  wire                IBusCachedPlugin_mmuBus_rsp_isIoAccess;
  wire                IBusCachedPlugin_mmuBus_rsp_isPaging;
  wire                IBusCachedPlugin_mmuBus_rsp_allowRead;
  wire                IBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire                IBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire                IBusCachedPlugin_mmuBus_rsp_exception;
  wire                IBusCachedPlugin_mmuBus_rsp_refilling;
  wire                IBusCachedPlugin_mmuBus_rsp_bypassTranslation;
  wire                IBusCachedPlugin_mmuBus_end;
  wire                IBusCachedPlugin_mmuBus_busy;
  reg                 DBusSimplePlugin_memoryExceptionPort_valid;
  reg        [3:0]    DBusSimplePlugin_memoryExceptionPort_payload_code;
  wire       [31:0]   DBusSimplePlugin_memoryExceptionPort_payload_badAddr;
  wire                decodeExceptionPort_valid;
  wire       [3:0]    decodeExceptionPort_payload_code;
  wire       [31:0]   decodeExceptionPort_payload_badAddr;
  wire                BranchPlugin_jumpInterface_valid;
  wire       [31:0]   BranchPlugin_jumpInterface_payload;
  wire                BranchPlugin_branchExceptionPort_valid;
  wire       [3:0]    BranchPlugin_branchExceptionPort_payload_code;
  wire       [31:0]   BranchPlugin_branchExceptionPort_payload_badAddr;
  wire       [31:0]   CsrPlugin_csrMapping_readDataSignal;
  wire       [31:0]   CsrPlugin_csrMapping_readDataInit;
  wire       [31:0]   CsrPlugin_csrMapping_writeDataSignal;
  wire                CsrPlugin_csrMapping_allowCsrSignal;
  wire                CsrPlugin_csrMapping_hazardFree;
  wire                CsrPlugin_inWfi /* verilator public */ ;
  reg                 CsrPlugin_thirdPartyWake;
  reg                 CsrPlugin_jumpInterface_valid;
  reg        [31:0]   CsrPlugin_jumpInterface_payload;
  wire                CsrPlugin_exceptionPendings_0;
  wire                CsrPlugin_exceptionPendings_1;
  wire                CsrPlugin_exceptionPendings_2;
  wire                CsrPlugin_exceptionPendings_3;
  wire                externalInterrupt;
  wire                contextSwitching;
  reg        [1:0]    CsrPlugin_privilege;
  reg                 CsrPlugin_forceMachineWire;
  reg                 CsrPlugin_selfException_valid;
  reg        [3:0]    CsrPlugin_selfException_payload_code;
  wire       [31:0]   CsrPlugin_selfException_payload_badAddr;
  reg                 CsrPlugin_allowInterrupts;
  reg                 CsrPlugin_allowException;
  reg                 CsrPlugin_allowEbreakException;
  reg                 IBusCachedPlugin_injectionPort_valid;
  reg                 IBusCachedPlugin_injectionPort_ready;
  wire       [31:0]   IBusCachedPlugin_injectionPort_payload;
  wire                IBusCachedPlugin_externalFlush;
  wire                IBusCachedPlugin_jump_pcLoad_valid;
  wire       [31:0]   IBusCachedPlugin_jump_pcLoad_payload;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload;
  wire                IBusCachedPlugin_fetchPc_output_valid;
  wire                IBusCachedPlugin_fetchPc_output_ready;
  wire       [31:0]   IBusCachedPlugin_fetchPc_output_payload;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pcReg /* verilator public */ ;
  reg                 IBusCachedPlugin_fetchPc_correction;
  reg                 IBusCachedPlugin_fetchPc_correctionReg;
  wire                IBusCachedPlugin_fetchPc_output_fire;
  wire                IBusCachedPlugin_fetchPc_corrected;
  reg                 IBusCachedPlugin_fetchPc_pcRegPropagate;
  reg                 IBusCachedPlugin_fetchPc_booted;
  reg                 IBusCachedPlugin_fetchPc_inc;
  wire                when_Fetcher_l131;
  wire                IBusCachedPlugin_fetchPc_output_fire_1;
  wire                when_Fetcher_l131_1;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pc;
  wire                IBusCachedPlugin_fetchPc_redo_valid;
  wire       [31:0]   IBusCachedPlugin_fetchPc_redo_payload;
  reg                 IBusCachedPlugin_fetchPc_flushed;
  wire                when_Fetcher_l158;
  reg                 IBusCachedPlugin_iBusRsp_redoFetch;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_0_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_1_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_2_halt;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire                IBusCachedPlugin_iBusRsp_flush;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  reg        [31:0]   _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 IBusCachedPlugin_iBusRsp_readyForError;
  wire                IBusCachedPlugin_iBusRsp_output_valid;
  wire                IBusCachedPlugin_iBusRsp_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_pc;
  wire                IBusCachedPlugin_iBusRsp_output_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  wire                IBusCachedPlugin_iBusRsp_output_payload_isRvc;
  wire                when_Fetcher_l240;
  wire                when_Fetcher_l320;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_0;
  wire                when_Fetcher_l329;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_1;
  wire                when_Fetcher_l329_1;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_2;
  wire                when_Fetcher_l329_2;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_3;
  wire                when_Fetcher_l329_3;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_4;
  wire                when_Fetcher_l329_4;
  wire                iBus_cmd_valid;
  wire                iBus_cmd_ready;
  reg        [31:0]   iBus_cmd_payload_address;
  wire       [2:0]    iBus_cmd_payload_size;
  wire                iBus_rsp_valid;
  wire       [31:0]   iBus_rsp_payload_data;
  wire                iBus_rsp_payload_error;
  wire       [31:0]   _zz_IBusCachedPlugin_rspCounter;
  reg        [31:0]   IBusCachedPlugin_rspCounter;
  wire                IBusCachedPlugin_s0_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s1_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s2_tightlyCoupledHit;
  wire                IBusCachedPlugin_rsp_iBusRspOutputHalt;
  wire                IBusCachedPlugin_rsp_issueDetected;
  reg                 IBusCachedPlugin_rsp_redoFetch;
  wire                when_IBusCachedPlugin_l239;
  wire                when_IBusCachedPlugin_l244;
  wire                when_IBusCachedPlugin_l250;
  wire                when_IBusCachedPlugin_l256;
  wire                when_IBusCachedPlugin_l267;
  wire                dBus_cmd_valid;
  wire                dBus_cmd_ready;
  wire                dBus_cmd_payload_wr;
  wire       [31:0]   dBus_cmd_payload_address;
  wire       [31:0]   dBus_cmd_payload_data;
  wire       [1:0]    dBus_cmd_payload_size;
  wire                dBus_rsp_ready;
  wire                dBus_rsp_error;
  wire       [31:0]   dBus_rsp_data;
  wire                _zz_dBus_cmd_valid;
  reg                 execute_DBusSimplePlugin_skipCmd;
  reg        [31:0]   _zz_dBus_cmd_payload_data;
  wire                when_DBusSimplePlugin_l426;
  reg        [3:0]    _zz_execute_DBusSimplePlugin_formalMask;
  wire       [3:0]    execute_DBusSimplePlugin_formalMask;
  wire                when_DBusSimplePlugin_l479;
  wire                when_DBusSimplePlugin_l486;
  wire                when_DBusSimplePlugin_l512;
  reg        [31:0]   writeBack_DBusSimplePlugin_rspShifted;
  wire       [1:0]    switch_Misc_l200;
  wire                _zz_writeBack_DBusSimplePlugin_rspFormated;
  reg        [31:0]   _zz_writeBack_DBusSimplePlugin_rspFormated_1;
  wire                _zz_writeBack_DBusSimplePlugin_rspFormated_2;
  reg        [31:0]   _zz_writeBack_DBusSimplePlugin_rspFormated_3;
  reg        [31:0]   writeBack_DBusSimplePlugin_rspFormated;
  wire                when_DBusSimplePlugin_l558;
  wire       [27:0]   _zz_decode_ENV_CTRL_2;
  wire                _zz_decode_ENV_CTRL_3;
  wire                _zz_decode_ENV_CTRL_4;
  wire                _zz_decode_ENV_CTRL_5;
  wire                _zz_decode_ENV_CTRL_6;
  wire       [1:0] _zz_decode_SRC1_CTRL_2;
  wire       [1:0] _zz_decode_ALU_CTRL_2;
  wire       [1:0] _zz_decode_SRC2_CTRL_2;
  wire       [1:0] _zz_decode_ALU_BITWISE_CTRL_2;
  wire       [1:0] _zz_decode_SHIFT_CTRL_2;
  wire       [1:0] _zz_decode_BRANCH_CTRL_2;
  wire       [1:0] _zz_decode_ENV_CTRL_7;
  wire                when_RegFilePlugin_l63;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress1;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress2;
  wire       [31:0]   decode_RegFilePlugin_rs1Data;
  wire       [31:0]   decode_RegFilePlugin_rs2Data;
  reg                 lastStageRegFileWrite_valid /* verilator public */ ;
  reg        [4:0]    lastStageRegFileWrite_payload_address /* verilator public */ ;
  reg        [31:0]   lastStageRegFileWrite_payload_data /* verilator public */ ;
  reg                 _zz_2;
  reg        [31:0]   execute_IntAluPlugin_bitwise;
  reg        [31:0]   _zz_execute_REGFILE_WRITE_DATA;
  reg        [31:0]   _zz_execute_SRC1;
  wire                _zz_execute_SRC2_1;
  reg        [19:0]   _zz_execute_SRC2_2;
  wire                _zz_execute_SRC2_3;
  reg        [19:0]   _zz_execute_SRC2_4;
  reg        [31:0]   _zz_execute_SRC2_5;
  reg        [31:0]   execute_SrcPlugin_addSub;
  wire                execute_SrcPlugin_less;
  reg                 execute_LightShifterPlugin_isActive;
  wire                execute_LightShifterPlugin_isShift;
  reg        [4:0]    execute_LightShifterPlugin_amplitudeReg;
  wire       [4:0]    execute_LightShifterPlugin_amplitude;
  wire       [31:0]   execute_LightShifterPlugin_shiftInput;
  wire                execute_LightShifterPlugin_done;
  wire                when_ShiftPlugins_l169;
  reg        [31:0]   _zz_execute_to_memory_REGFILE_WRITE_DATA_1;
  wire                when_ShiftPlugins_l175;
  wire                when_ShiftPlugins_l184;
  reg                 HazardSimplePlugin_src0Hazard;
  reg                 HazardSimplePlugin_src1Hazard;
  wire                HazardSimplePlugin_writeBackWrites_valid;
  wire       [4:0]    HazardSimplePlugin_writeBackWrites_payload_address;
  wire       [31:0]   HazardSimplePlugin_writeBackWrites_payload_data;
  reg                 HazardSimplePlugin_writeBackBuffer_valid;
  reg        [4:0]    HazardSimplePlugin_writeBackBuffer_payload_address;
  reg        [31:0]   HazardSimplePlugin_writeBackBuffer_payload_data;
  wire                HazardSimplePlugin_addr0Match;
  wire                HazardSimplePlugin_addr1Match;
  wire                when_HazardSimplePlugin_l59;
  wire                when_HazardSimplePlugin_l62;
  wire                when_HazardSimplePlugin_l57;
  wire                when_HazardSimplePlugin_l58;
  wire                when_HazardSimplePlugin_l59_1;
  wire                when_HazardSimplePlugin_l62_1;
  wire                when_HazardSimplePlugin_l57_1;
  wire                when_HazardSimplePlugin_l58_1;
  wire                when_HazardSimplePlugin_l59_2;
  wire                when_HazardSimplePlugin_l62_2;
  wire                when_HazardSimplePlugin_l57_2;
  wire                when_HazardSimplePlugin_l58_2;
  wire                when_HazardSimplePlugin_l105;
  wire                when_HazardSimplePlugin_l108;
  wire                when_HazardSimplePlugin_l113;
  wire                execute_BranchPlugin_eq;
  wire       [2:0]    switch_Misc_l200_1;
  reg                 _zz_execute_BRANCH_DO;
  reg                 _zz_execute_BRANCH_DO_1;
  wire       [31:0]   execute_BranchPlugin_branch_src1;
  wire                _zz_execute_BranchPlugin_branch_src2;
  reg        [10:0]   _zz_execute_BranchPlugin_branch_src2_1;
  wire                _zz_execute_BranchPlugin_branch_src2_2;
  reg        [19:0]   _zz_execute_BranchPlugin_branch_src2_3;
  wire                _zz_execute_BranchPlugin_branch_src2_4;
  reg        [18:0]   _zz_execute_BranchPlugin_branch_src2_5;
  reg        [31:0]   _zz_execute_BranchPlugin_branch_src2_6;
  wire       [31:0]   execute_BranchPlugin_branch_src2;
  wire       [31:0]   execute_BranchPlugin_branchAdder;
  wire       [1:0]    CsrPlugin_misa_base;
  wire       [25:0]   CsrPlugin_misa_extensions;
  reg        [1:0]    CsrPlugin_mtvec_mode;
  reg        [29:0]   CsrPlugin_mtvec_base;
  reg        [31:0]   CsrPlugin_mepc;
  reg                 CsrPlugin_mstatus_MIE;
  reg                 CsrPlugin_mstatus_MPIE;
  reg        [1:0]    CsrPlugin_mstatus_MPP;
  reg                 CsrPlugin_mip_MEIP;
  reg                 CsrPlugin_mip_MTIP;
  reg                 CsrPlugin_mip_MSIP;
  reg                 CsrPlugin_mie_MEIE;
  reg                 CsrPlugin_mie_MTIE;
  reg                 CsrPlugin_mie_MSIE;
  reg                 CsrPlugin_mcause_interrupt;
  reg        [3:0]    CsrPlugin_mcause_exceptionCode;
  reg        [31:0]   CsrPlugin_mtval;
  reg        [63:0]   CsrPlugin_mcycle = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  reg        [63:0]   CsrPlugin_minstret = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire                _zz_when_CsrPlugin_l952;
  wire                _zz_when_CsrPlugin_l952_1;
  wire                _zz_when_CsrPlugin_l952_2;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  reg        [3:0]    CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  reg        [31:0]   CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
  wire       [1:0]    _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  wire                _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire       [1:0]    _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_2;
  wire                _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3;
  wire                when_CsrPlugin_l909;
  wire                when_CsrPlugin_l909_1;
  wire                when_CsrPlugin_l909_2;
  wire                when_CsrPlugin_l909_3;
  wire                when_CsrPlugin_l922;
  reg                 CsrPlugin_interrupt_valid;
  reg        [3:0]    CsrPlugin_interrupt_code /* verilator public */ ;
  reg        [1:0]    CsrPlugin_interrupt_targetPrivilege;
  wire                when_CsrPlugin_l946;
  wire                when_CsrPlugin_l952;
  wire                when_CsrPlugin_l952_1;
  wire                when_CsrPlugin_l952_2;
  wire                CsrPlugin_exception;
  wire                CsrPlugin_lastStageWasWfi;
  reg                 CsrPlugin_pipelineLiberator_pcValids_0;
  reg                 CsrPlugin_pipelineLiberator_pcValids_1;
  reg                 CsrPlugin_pipelineLiberator_pcValids_2;
  wire                CsrPlugin_pipelineLiberator_active;
  wire                when_CsrPlugin_l980;
  wire                when_CsrPlugin_l980_1;
  wire                when_CsrPlugin_l980_2;
  wire                when_CsrPlugin_l985;
  reg                 CsrPlugin_pipelineLiberator_done;
  wire                when_CsrPlugin_l991;
  wire                CsrPlugin_interruptJump /* verilator public */ ;
  reg                 CsrPlugin_hadException /* verilator public */ ;
  reg        [1:0]    CsrPlugin_targetPrivilege;
  reg        [3:0]    CsrPlugin_trapCause;
  reg        [1:0]    CsrPlugin_xtvec_mode;
  reg        [29:0]   CsrPlugin_xtvec_base;
  wire                when_CsrPlugin_l1019;
  wire                when_CsrPlugin_l1064;
  wire       [1:0]    switch_CsrPlugin_l1068;
  reg                 execute_CsrPlugin_wfiWake;
  wire                when_CsrPlugin_l1116;
  wire                execute_CsrPlugin_blockedBySideEffects;
  reg                 execute_CsrPlugin_illegalAccess;
  reg                 execute_CsrPlugin_illegalInstruction;
  wire                when_CsrPlugin_l1136;
  wire                when_CsrPlugin_l1137;
  wire                when_CsrPlugin_l1144;
  reg                 execute_CsrPlugin_writeInstruction;
  reg                 execute_CsrPlugin_readInstruction;
  wire                execute_CsrPlugin_writeEnable;
  wire                execute_CsrPlugin_readEnable;
  wire       [31:0]   execute_CsrPlugin_readToWriteData;
  wire                switch_Misc_l200_2;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_writeDataSignal;
  wire                when_CsrPlugin_l1176;
  wire                when_CsrPlugin_l1180;
  wire       [11:0]   execute_CsrPlugin_csrAddress;
  reg        [31:0]   externalInterruptArray_regNext;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_1;
  reg                 DebugPlugin_firstCycle;
  reg                 DebugPlugin_secondCycle;
  reg                 DebugPlugin_resetIt;
  reg                 DebugPlugin_haltIt;
  reg                 DebugPlugin_stepIt;
  reg                 DebugPlugin_isPipBusy;
  reg                 DebugPlugin_godmode;
  wire                when_DebugPlugin_l225;
  reg                 DebugPlugin_haltedByBreak;
  reg                 DebugPlugin_debugUsed /* verilator public */ ;
  reg                 DebugPlugin_disableEbreak;
  wire                DebugPlugin_allowEBreak;
  reg        [31:0]   DebugPlugin_busReadDataReg;
  reg                 _zz_when_DebugPlugin_l244;
  wire                when_DebugPlugin_l244;
  wire       [5:0]    switch_DebugPlugin_l256;
  wire                when_DebugPlugin_l260;
  wire                when_DebugPlugin_l260_1;
  wire                when_DebugPlugin_l261;
  wire                when_DebugPlugin_l261_1;
  wire                when_DebugPlugin_l262;
  wire                when_DebugPlugin_l263;
  wire                when_DebugPlugin_l264;
  wire                when_DebugPlugin_l264_1;
  wire                when_DebugPlugin_l284;
  wire                when_DebugPlugin_l287;
  wire                when_DebugPlugin_l300;
  reg                 DebugPlugin_resetIt_regNext;
  wire                when_DebugPlugin_l316;
  wire                when_Pipeline_l124;
  reg        [31:0]   decode_to_execute_PC;
  wire                when_Pipeline_l124_1;
  reg        [31:0]   execute_to_memory_PC;
  wire                when_Pipeline_l124_2;
  reg        [31:0]   memory_to_writeBack_PC;
  wire                when_Pipeline_l124_3;
  reg        [31:0]   decode_to_execute_INSTRUCTION;
  wire                when_Pipeline_l124_4;
  reg        [31:0]   execute_to_memory_INSTRUCTION;
  wire                when_Pipeline_l124_5;
  reg        [31:0]   memory_to_writeBack_INSTRUCTION;
  wire                when_Pipeline_l124_6;
  reg        [31:0]   decode_to_execute_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_7;
  reg        [31:0]   execute_to_memory_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_8;
  reg        [31:0]   memory_to_writeBack_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_9;
  reg        [1:0] decode_to_execute_SRC1_CTRL;
  wire                when_Pipeline_l124_10;
  reg                 decode_to_execute_SRC_USE_SUB_LESS;
  wire                when_Pipeline_l124_11;
  reg                 decode_to_execute_MEMORY_ENABLE;
  wire                when_Pipeline_l124_12;
  reg                 execute_to_memory_MEMORY_ENABLE;
  wire                when_Pipeline_l124_13;
  reg                 memory_to_writeBack_MEMORY_ENABLE;
  wire                when_Pipeline_l124_14;
  reg        [1:0] decode_to_execute_ALU_CTRL;
  wire                when_Pipeline_l124_15;
  reg        [1:0] decode_to_execute_SRC2_CTRL;
  wire                when_Pipeline_l124_16;
  reg                 decode_to_execute_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_17;
  reg                 execute_to_memory_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_18;
  reg                 memory_to_writeBack_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_19;
  reg                 decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  wire                when_Pipeline_l124_20;
  reg                 decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_21;
  reg                 execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_22;
  reg                 decode_to_execute_MEMORY_STORE;
  wire                when_Pipeline_l124_23;
  reg                 execute_to_memory_MEMORY_STORE;
  wire                when_Pipeline_l124_24;
  reg                 memory_to_writeBack_MEMORY_STORE;
  wire                when_Pipeline_l124_25;
  reg                 decode_to_execute_SRC_LESS_UNSIGNED;
  wire                when_Pipeline_l124_26;
  reg        [1:0] decode_to_execute_ALU_BITWISE_CTRL;
  wire                when_Pipeline_l124_27;
  reg        [1:0] decode_to_execute_SHIFT_CTRL;
  wire                when_Pipeline_l124_28;
  reg        [1:0] decode_to_execute_BRANCH_CTRL;
  wire                when_Pipeline_l124_29;
  reg                 decode_to_execute_IS_CSR;
  wire                when_Pipeline_l124_30;
  reg        [1:0] decode_to_execute_ENV_CTRL;
  wire                when_Pipeline_l124_31;
  reg        [1:0] execute_to_memory_ENV_CTRL;
  wire                when_Pipeline_l124_32;
  reg        [1:0] memory_to_writeBack_ENV_CTRL;
  wire                when_Pipeline_l124_33;
  reg        [31:0]   decode_to_execute_RS1;
  wire                when_Pipeline_l124_34;
  reg        [31:0]   decode_to_execute_RS2;
  wire                when_Pipeline_l124_35;
  reg                 decode_to_execute_SRC2_FORCE_ZERO;
  wire                when_Pipeline_l124_36;
  reg                 decode_to_execute_CSR_WRITE_OPCODE;
  wire                when_Pipeline_l124_37;
  reg                 decode_to_execute_CSR_READ_OPCODE;
  wire                when_Pipeline_l124_38;
  reg                 decode_to_execute_DO_EBREAK;
  wire                when_Pipeline_l124_39;
  reg                 execute_to_memory_ALIGNEMENT_FAULT;
  wire                when_Pipeline_l124_40;
  reg        [1:0]    execute_to_memory_MEMORY_ADDRESS_LOW;
  wire                when_Pipeline_l124_41;
  reg        [1:0]    memory_to_writeBack_MEMORY_ADDRESS_LOW;
  wire                when_Pipeline_l124_42;
  reg        [31:0]   execute_to_memory_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_43;
  reg        [31:0]   memory_to_writeBack_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_44;
  reg                 execute_to_memory_BRANCH_DO;
  wire                when_Pipeline_l124_45;
  reg        [31:0]   execute_to_memory_BRANCH_CALC;
  wire                when_Pipeline_l124_46;
  reg        [31:0]   memory_to_writeBack_MEMORY_READ_DATA;
  wire                when_Pipeline_l151;
  wire                when_Pipeline_l154;
  wire                when_Pipeline_l151_1;
  wire                when_Pipeline_l154_1;
  wire                when_Pipeline_l151_2;
  wire                when_Pipeline_l154_2;
  reg        [2:0]    switch_Fetcher_l362;
  wire                when_Fetcher_l378;
  wire                when_CsrPlugin_l1264;
  reg                 execute_CsrPlugin_csr_768;
  wire                when_CsrPlugin_l1264_1;
  reg                 execute_CsrPlugin_csr_836;
  wire                when_CsrPlugin_l1264_2;
  reg                 execute_CsrPlugin_csr_772;
  wire                when_CsrPlugin_l1264_3;
  reg                 execute_CsrPlugin_csr_773;
  wire                when_CsrPlugin_l1264_4;
  reg                 execute_CsrPlugin_csr_833;
  wire                when_CsrPlugin_l1264_5;
  reg                 execute_CsrPlugin_csr_834;
  wire                when_CsrPlugin_l1264_6;
  reg                 execute_CsrPlugin_csr_835;
  wire                when_CsrPlugin_l1264_7;
  reg                 execute_CsrPlugin_csr_3008;
  wire                when_CsrPlugin_l1264_8;
  reg                 execute_CsrPlugin_csr_4032;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_2;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_3;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_4;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_5;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_6;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_7;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_8;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_9;
  wire                when_CsrPlugin_l1297;
  wire                when_CsrPlugin_l1302;
  reg        [2:0]    _zz_iBusWishbone_ADR;
  wire                when_InstructionCache_l239;
  reg                 _zz_iBus_rsp_valid;
  reg        [31:0]   iBusWishbone_DAT_MISO_regNext;
  wire                dBus_cmd_halfPipe_valid;
  wire                dBus_cmd_halfPipe_ready;
  wire                dBus_cmd_halfPipe_payload_wr;
  wire       [31:0]   dBus_cmd_halfPipe_payload_address;
  wire       [31:0]   dBus_cmd_halfPipe_payload_data;
  wire       [1:0]    dBus_cmd_halfPipe_payload_size;
  reg                 dBus_cmd_rValid;
  wire                dBus_cmd_halfPipe_fire;
  reg                 dBus_cmd_rData_wr;
  reg        [31:0]   dBus_cmd_rData_address;
  reg        [31:0]   dBus_cmd_rData_data;
  reg        [1:0]    dBus_cmd_rData_size;
  reg        [3:0]    _zz_dBusWishbone_SEL;
  wire                when_DBusSimplePlugin_l189;
  
  reg [39:0] _zz_memory_to_writeBack_ENV_CTRL_string;
  reg [39:0] _zz_memory_to_writeBack_ENV_CTRL_1_string;
  reg [39:0] _zz_execute_to_memory_ENV_CTRL_string;
  reg [39:0] _zz_execute_to_memory_ENV_CTRL_1_string;
  reg [39:0] decode_ENV_CTRL_string;
  reg [39:0] _zz_decode_ENV_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ENV_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ENV_CTRL_1_string;
  reg [31:0] decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_1_string;
  reg [71:0] decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_1_string;
  reg [39:0] decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string;
  reg [23:0] decode_SRC2_CTRL_string;
  reg [23:0] _zz_decode_SRC2_CTRL_string;
  reg [23:0] _zz_decode_to_execute_SRC2_CTRL_string;
  reg [23:0] _zz_decode_to_execute_SRC2_CTRL_1_string;
  reg [63:0] decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_1_string;
  reg [95:0] decode_SRC1_CTRL_string;
  reg [95:0] _zz_decode_SRC1_CTRL_string;
  reg [95:0] _zz_decode_to_execute_SRC1_CTRL_string;
  reg [95:0] _zz_decode_to_execute_SRC1_CTRL_1_string;
  reg [39:0] memory_ENV_CTRL_string;
  reg [39:0] _zz_memory_ENV_CTRL_string;
  reg [39:0] execute_ENV_CTRL_string;
  reg [39:0] _zz_execute_ENV_CTRL_string;
  reg [39:0] writeBack_ENV_CTRL_string;
  reg [39:0] _zz_writeBack_ENV_CTRL_string;
  reg [31:0] execute_BRANCH_CTRL_string;
  reg [31:0] _zz_execute_BRANCH_CTRL_string;
  reg [71:0] execute_SHIFT_CTRL_string;
  reg [71:0] _zz_execute_SHIFT_CTRL_string;
  reg [23:0] execute_SRC2_CTRL_string;
  reg [23:0] _zz_execute_SRC2_CTRL_string;
  reg [95:0] execute_SRC1_CTRL_string;
  reg [95:0] _zz_execute_SRC1_CTRL_string;
  reg [63:0] execute_ALU_CTRL_string;
  reg [63:0] _zz_execute_ALU_CTRL_string;
  reg [39:0] execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_ENV_CTRL_1_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_1_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_1_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_1_string;
  reg [23:0] _zz_decode_SRC2_CTRL_1_string;
  reg [63:0] _zz_decode_ALU_CTRL_1_string;
  reg [95:0] _zz_decode_SRC1_CTRL_1_string;
  reg [95:0] _zz_decode_SRC1_CTRL_2_string;
  reg [63:0] _zz_decode_ALU_CTRL_2_string;
  reg [23:0] _zz_decode_SRC2_CTRL_2_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_2_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_2_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_2_string;
  reg [39:0] _zz_decode_ENV_CTRL_7_string;
  reg [95:0] decode_to_execute_SRC1_CTRL_string;
  reg [63:0] decode_to_execute_ALU_CTRL_string;
  reg [23:0] decode_to_execute_SRC2_CTRL_string;
  reg [39:0] decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [71:0] decode_to_execute_SHIFT_CTRL_string;
  reg [31:0] decode_to_execute_BRANCH_CTRL_string;
  reg [39:0] decode_to_execute_ENV_CTRL_string;
  reg [39:0] execute_to_memory_ENV_CTRL_string;
  reg [39:0] memory_to_writeBack_ENV_CTRL_string;
  

  (* ram_style = "block" *) reg [31:0] RegFilePlugin_regFile [0:31] /* verilator public */ ;

  assign _zz_when = ({decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid} != 2'b00);
  assign _zz_when_1 = ({BranchPlugin_branchExceptionPort_valid,DBusSimplePlugin_memoryExceptionPort_valid} != 2'b00);
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_1 = (_zz_IBusCachedPlugin_jump_pcLoad_payload & (~ _zz_IBusCachedPlugin_jump_pcLoad_payload_2));
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_2 = (_zz_IBusCachedPlugin_jump_pcLoad_payload - 2'b01);
  assign _zz_IBusCachedPlugin_fetchPc_pc_1 = {IBusCachedPlugin_fetchPc_inc,2'b00};
  assign _zz_IBusCachedPlugin_fetchPc_pc = {29'd0, _zz_IBusCachedPlugin_fetchPc_pc_1};
  assign _zz_DBusSimplePlugin_memoryExceptionPort_payload_code = (memory_MEMORY_STORE ? 3'b110 : 3'b100);
  assign _zz__zz_execute_REGFILE_WRITE_DATA = execute_SRC_LESS;
  assign _zz__zz_execute_SRC1 = 3'b100;
  assign _zz__zz_execute_SRC1_1 = execute_INSTRUCTION[19 : 15];
  assign _zz__zz_execute_SRC2_3 = {execute_INSTRUCTION[31 : 25],execute_INSTRUCTION[11 : 7]};
  assign _zz_execute_SrcPlugin_addSub = ($signed(_zz_execute_SrcPlugin_addSub_1) + $signed(_zz_execute_SrcPlugin_addSub_4));
  assign _zz_execute_SrcPlugin_addSub_1 = ($signed(_zz_execute_SrcPlugin_addSub_2) + $signed(_zz_execute_SrcPlugin_addSub_3));
  assign _zz_execute_SrcPlugin_addSub_2 = execute_SRC1;
  assign _zz_execute_SrcPlugin_addSub_3 = (execute_SRC_USE_SUB_LESS ? (~ execute_SRC2) : execute_SRC2);
  assign _zz_execute_SrcPlugin_addSub_4 = (execute_SRC_USE_SUB_LESS ? _zz_execute_SrcPlugin_addSub_5 : _zz_execute_SrcPlugin_addSub_6);
  assign _zz_execute_SrcPlugin_addSub_5 = 32'h00000001;
  assign _zz_execute_SrcPlugin_addSub_6 = 32'h0;
  assign _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1 = (_zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1_1 >>> 1);
  assign _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1_1 = {((execute_SHIFT_CTRL == 2'b11) && execute_LightShifterPlugin_shiftInput[31]),execute_LightShifterPlugin_shiftInput};
  assign _zz__zz_execute_BranchPlugin_branch_src2 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]};
  assign _zz__zz_execute_BranchPlugin_branch_src2_4 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]};
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code & (~ _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1));
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code - 2'b01);
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_2 & (~ _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3_1));
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_2 - 2'b01);
  assign _zz_iBusWishbone_ADR_1 = (iBus_cmd_payload_address >>> 5);
  assign _zz_decode_RegFilePlugin_rs1Data = 1'b1;
  assign _zz_decode_RegFilePlugin_rs2Data = 1'b1;
  assign _zz_decode_LEGAL_INSTRUCTION = 32'h0000107f;
  assign _zz_decode_LEGAL_INSTRUCTION_1 = (decode_INSTRUCTION & 32'h0000207f);
  assign _zz_decode_LEGAL_INSTRUCTION_2 = 32'h00002073;
  assign _zz_decode_LEGAL_INSTRUCTION_3 = ((decode_INSTRUCTION & 32'h0000407f) == 32'h00004063);
  assign _zz_decode_LEGAL_INSTRUCTION_4 = ((decode_INSTRUCTION & 32'h0000207f) == 32'h00002013);
  assign _zz_decode_LEGAL_INSTRUCTION_5 = {((decode_INSTRUCTION & 32'h0000603f) == 32'h00000023),{((decode_INSTRUCTION & 32'h0000207f) == 32'h00000003),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_6) == 32'h00000003),{(_zz_decode_LEGAL_INSTRUCTION_7 == _zz_decode_LEGAL_INSTRUCTION_8),{_zz_decode_LEGAL_INSTRUCTION_9,{_zz_decode_LEGAL_INSTRUCTION_10,_zz_decode_LEGAL_INSTRUCTION_11}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_6 = 32'h0000505f;
  assign _zz_decode_LEGAL_INSTRUCTION_7 = (decode_INSTRUCTION & 32'h0000707b);
  assign _zz_decode_LEGAL_INSTRUCTION_8 = 32'h00000063;
  assign _zz_decode_LEGAL_INSTRUCTION_9 = ((decode_INSTRUCTION & 32'h0000607f) == 32'h0000000f);
  assign _zz_decode_LEGAL_INSTRUCTION_10 = ((decode_INSTRUCTION & 32'hfe00007f) == 32'h00000033);
  assign _zz_decode_LEGAL_INSTRUCTION_11 = {((decode_INSTRUCTION & 32'hbc00707f) == 32'h00005013),{((decode_INSTRUCTION & 32'hfc00307f) == 32'h00001013),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_12) == 32'h00005033),{(_zz_decode_LEGAL_INSTRUCTION_13 == _zz_decode_LEGAL_INSTRUCTION_14),{_zz_decode_LEGAL_INSTRUCTION_15,{_zz_decode_LEGAL_INSTRUCTION_16,_zz_decode_LEGAL_INSTRUCTION_17}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_12 = 32'hbe00707f;
  assign _zz_decode_LEGAL_INSTRUCTION_13 = (decode_INSTRUCTION & 32'hbe00707f);
  assign _zz_decode_LEGAL_INSTRUCTION_14 = 32'h00000033;
  assign _zz_decode_LEGAL_INSTRUCTION_15 = ((decode_INSTRUCTION & 32'hdfffffff) == 32'h10200073);
  assign _zz_decode_LEGAL_INSTRUCTION_16 = ((decode_INSTRUCTION & 32'hffefffff) == 32'h00000073);
  assign _zz_decode_LEGAL_INSTRUCTION_17 = ((decode_INSTRUCTION & 32'hffffffff) == 32'h10500073);
  assign _zz__zz_decode_ENV_CTRL_2 = 32'h10103050;
  assign _zz__zz_decode_ENV_CTRL_2_1 = (decode_INSTRUCTION & 32'h10103050);
  assign _zz__zz_decode_ENV_CTRL_2_2 = 32'h00000050;
  assign _zz__zz_decode_ENV_CTRL_2_3 = ((decode_INSTRUCTION & 32'h10403050) == 32'h10000050);
  assign _zz__zz_decode_ENV_CTRL_2_4 = {(_zz__zz_decode_ENV_CTRL_2_5 == _zz__zz_decode_ENV_CTRL_2_6),(_zz__zz_decode_ENV_CTRL_2_7 == _zz__zz_decode_ENV_CTRL_2_8)};
  assign _zz__zz_decode_ENV_CTRL_2_9 = 2'b00;
  assign _zz__zz_decode_ENV_CTRL_2_10 = ({_zz_decode_ENV_CTRL_6,_zz__zz_decode_ENV_CTRL_2_11} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_12 = (_zz__zz_decode_ENV_CTRL_2_13 != 1'b0);
  assign _zz__zz_decode_ENV_CTRL_2_14 = {(_zz__zz_decode_ENV_CTRL_2_15 != _zz__zz_decode_ENV_CTRL_2_17),{_zz__zz_decode_ENV_CTRL_2_18,{_zz__zz_decode_ENV_CTRL_2_21,_zz__zz_decode_ENV_CTRL_2_26}}};
  assign _zz__zz_decode_ENV_CTRL_2_5 = (decode_INSTRUCTION & 32'h00001050);
  assign _zz__zz_decode_ENV_CTRL_2_6 = 32'h00001050;
  assign _zz__zz_decode_ENV_CTRL_2_7 = (decode_INSTRUCTION & 32'h00002050);
  assign _zz__zz_decode_ENV_CTRL_2_8 = 32'h00002050;
  assign _zz__zz_decode_ENV_CTRL_2_11 = ((decode_INSTRUCTION & 32'h0000001c) == 32'h00000004);
  assign _zz__zz_decode_ENV_CTRL_2_13 = ((decode_INSTRUCTION & 32'h00000058) == 32'h00000040);
  assign _zz__zz_decode_ENV_CTRL_2_15 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_16) == 32'h00005010);
  assign _zz__zz_decode_ENV_CTRL_2_17 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_18 = ({_zz__zz_decode_ENV_CTRL_2_19,_zz__zz_decode_ENV_CTRL_2_20} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_21 = ({_zz__zz_decode_ENV_CTRL_2_22,_zz__zz_decode_ENV_CTRL_2_24} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_26 = {(_zz__zz_decode_ENV_CTRL_2_27 != _zz__zz_decode_ENV_CTRL_2_29),{_zz__zz_decode_ENV_CTRL_2_30,{_zz__zz_decode_ENV_CTRL_2_33,_zz__zz_decode_ENV_CTRL_2_38}}};
  assign _zz__zz_decode_ENV_CTRL_2_16 = 32'h00007054;
  assign _zz__zz_decode_ENV_CTRL_2_19 = ((decode_INSTRUCTION & 32'h40003054) == 32'h40001010);
  assign _zz__zz_decode_ENV_CTRL_2_20 = ((decode_INSTRUCTION & 32'h00007054) == 32'h00001010);
  assign _zz__zz_decode_ENV_CTRL_2_22 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_23) == 32'h00000024);
  assign _zz__zz_decode_ENV_CTRL_2_24 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_25) == 32'h00001010);
  assign _zz__zz_decode_ENV_CTRL_2_27 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_28) == 32'h00001000);
  assign _zz__zz_decode_ENV_CTRL_2_29 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_30 = ((_zz__zz_decode_ENV_CTRL_2_31 == _zz__zz_decode_ENV_CTRL_2_32) != 1'b0);
  assign _zz__zz_decode_ENV_CTRL_2_33 = ({_zz__zz_decode_ENV_CTRL_2_34,_zz__zz_decode_ENV_CTRL_2_36} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_38 = {(_zz__zz_decode_ENV_CTRL_2_39 != _zz__zz_decode_ENV_CTRL_2_44),{_zz__zz_decode_ENV_CTRL_2_45,{_zz__zz_decode_ENV_CTRL_2_51,_zz__zz_decode_ENV_CTRL_2_53}}};
  assign _zz__zz_decode_ENV_CTRL_2_23 = 32'h00000064;
  assign _zz__zz_decode_ENV_CTRL_2_25 = 32'h00003054;
  assign _zz__zz_decode_ENV_CTRL_2_28 = 32'h00001000;
  assign _zz__zz_decode_ENV_CTRL_2_31 = (decode_INSTRUCTION & 32'h00003000);
  assign _zz__zz_decode_ENV_CTRL_2_32 = 32'h00002000;
  assign _zz__zz_decode_ENV_CTRL_2_34 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_35) == 32'h00002000);
  assign _zz__zz_decode_ENV_CTRL_2_36 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_37) == 32'h00001000);
  assign _zz__zz_decode_ENV_CTRL_2_39 = {(_zz__zz_decode_ENV_CTRL_2_40 == _zz__zz_decode_ENV_CTRL_2_41),(_zz__zz_decode_ENV_CTRL_2_42 == _zz__zz_decode_ENV_CTRL_2_43)};
  assign _zz__zz_decode_ENV_CTRL_2_44 = 2'b00;
  assign _zz__zz_decode_ENV_CTRL_2_45 = ({_zz__zz_decode_ENV_CTRL_2_46,{_zz__zz_decode_ENV_CTRL_2_47,_zz__zz_decode_ENV_CTRL_2_49}} != 3'b000);
  assign _zz__zz_decode_ENV_CTRL_2_51 = (_zz__zz_decode_ENV_CTRL_2_52 != 1'b0);
  assign _zz__zz_decode_ENV_CTRL_2_53 = {(_zz__zz_decode_ENV_CTRL_2_54 != _zz__zz_decode_ENV_CTRL_2_56),{_zz__zz_decode_ENV_CTRL_2_57,{_zz__zz_decode_ENV_CTRL_2_58,_zz__zz_decode_ENV_CTRL_2_69}}};
  assign _zz__zz_decode_ENV_CTRL_2_35 = 32'h00002010;
  assign _zz__zz_decode_ENV_CTRL_2_37 = 32'h00005000;
  assign _zz__zz_decode_ENV_CTRL_2_40 = (decode_INSTRUCTION & 32'h00000034);
  assign _zz__zz_decode_ENV_CTRL_2_41 = 32'h00000020;
  assign _zz__zz_decode_ENV_CTRL_2_42 = (decode_INSTRUCTION & 32'h00000064);
  assign _zz__zz_decode_ENV_CTRL_2_43 = 32'h00000020;
  assign _zz__zz_decode_ENV_CTRL_2_46 = ((decode_INSTRUCTION & 32'h00000050) == 32'h00000040);
  assign _zz__zz_decode_ENV_CTRL_2_47 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_48) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_49 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_50) == 32'h00000040);
  assign _zz__zz_decode_ENV_CTRL_2_52 = ((decode_INSTRUCTION & 32'h00000020) == 32'h00000020);
  assign _zz__zz_decode_ENV_CTRL_2_54 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_55) == 32'h00000010);
  assign _zz__zz_decode_ENV_CTRL_2_56 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_57 = (_zz_decode_ENV_CTRL_5 != 1'b0);
  assign _zz__zz_decode_ENV_CTRL_2_58 = ({_zz__zz_decode_ENV_CTRL_2_59,_zz__zz_decode_ENV_CTRL_2_60} != 6'h0);
  assign _zz__zz_decode_ENV_CTRL_2_69 = {(_zz__zz_decode_ENV_CTRL_2_70 != _zz__zz_decode_ENV_CTRL_2_73),{_zz__zz_decode_ENV_CTRL_2_74,{_zz__zz_decode_ENV_CTRL_2_77,_zz__zz_decode_ENV_CTRL_2_84}}};
  assign _zz__zz_decode_ENV_CTRL_2_48 = 32'h00000038;
  assign _zz__zz_decode_ENV_CTRL_2_50 = 32'h00103040;
  assign _zz__zz_decode_ENV_CTRL_2_55 = 32'h00000010;
  assign _zz__zz_decode_ENV_CTRL_2_59 = _zz_decode_ENV_CTRL_6;
  assign _zz__zz_decode_ENV_CTRL_2_60 = {(_zz__zz_decode_ENV_CTRL_2_61 == _zz__zz_decode_ENV_CTRL_2_62),{_zz__zz_decode_ENV_CTRL_2_63,{_zz__zz_decode_ENV_CTRL_2_65,_zz__zz_decode_ENV_CTRL_2_66}}};
  assign _zz__zz_decode_ENV_CTRL_2_70 = {_zz_decode_ENV_CTRL_4,(_zz__zz_decode_ENV_CTRL_2_71 == _zz__zz_decode_ENV_CTRL_2_72)};
  assign _zz__zz_decode_ENV_CTRL_2_73 = 2'b00;
  assign _zz__zz_decode_ENV_CTRL_2_74 = ({_zz_decode_ENV_CTRL_4,_zz__zz_decode_ENV_CTRL_2_75} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_77 = ({_zz__zz_decode_ENV_CTRL_2_78,_zz__zz_decode_ENV_CTRL_2_81} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_84 = {(_zz__zz_decode_ENV_CTRL_2_85 != _zz__zz_decode_ENV_CTRL_2_88),{_zz__zz_decode_ENV_CTRL_2_89,{_zz__zz_decode_ENV_CTRL_2_97,_zz__zz_decode_ENV_CTRL_2_101}}};
  assign _zz__zz_decode_ENV_CTRL_2_61 = (decode_INSTRUCTION & 32'h00001010);
  assign _zz__zz_decode_ENV_CTRL_2_62 = 32'h00001010;
  assign _zz__zz_decode_ENV_CTRL_2_63 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_64) == 32'h00002010);
  assign _zz__zz_decode_ENV_CTRL_2_65 = _zz_decode_ENV_CTRL_5;
  assign _zz__zz_decode_ENV_CTRL_2_66 = {_zz__zz_decode_ENV_CTRL_2_67,_zz__zz_decode_ENV_CTRL_2_68};
  assign _zz__zz_decode_ENV_CTRL_2_71 = (decode_INSTRUCTION & 32'h00000070);
  assign _zz__zz_decode_ENV_CTRL_2_72 = 32'h00000020;
  assign _zz__zz_decode_ENV_CTRL_2_75 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_76) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_78 = (_zz__zz_decode_ENV_CTRL_2_79 == _zz__zz_decode_ENV_CTRL_2_80);
  assign _zz__zz_decode_ENV_CTRL_2_81 = (_zz__zz_decode_ENV_CTRL_2_82 == _zz__zz_decode_ENV_CTRL_2_83);
  assign _zz__zz_decode_ENV_CTRL_2_85 = (_zz__zz_decode_ENV_CTRL_2_86 == _zz__zz_decode_ENV_CTRL_2_87);
  assign _zz__zz_decode_ENV_CTRL_2_88 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_89 = ({_zz__zz_decode_ENV_CTRL_2_90,_zz__zz_decode_ENV_CTRL_2_92} != 4'b0000);
  assign _zz__zz_decode_ENV_CTRL_2_97 = (_zz__zz_decode_ENV_CTRL_2_98 != _zz__zz_decode_ENV_CTRL_2_100);
  assign _zz__zz_decode_ENV_CTRL_2_101 = {_zz__zz_decode_ENV_CTRL_2_102,{_zz__zz_decode_ENV_CTRL_2_108,_zz__zz_decode_ENV_CTRL_2_112}};
  assign _zz__zz_decode_ENV_CTRL_2_64 = 32'h00002010;
  assign _zz__zz_decode_ENV_CTRL_2_67 = ((decode_INSTRUCTION & 32'h0000000c) == 32'h00000004);
  assign _zz__zz_decode_ENV_CTRL_2_68 = ((decode_INSTRUCTION & 32'h00000028) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_76 = 32'h00000020;
  assign _zz__zz_decode_ENV_CTRL_2_79 = (decode_INSTRUCTION & 32'h00006014);
  assign _zz__zz_decode_ENV_CTRL_2_80 = 32'h00006010;
  assign _zz__zz_decode_ENV_CTRL_2_82 = (decode_INSTRUCTION & 32'h00005014);
  assign _zz__zz_decode_ENV_CTRL_2_83 = 32'h00004010;
  assign _zz__zz_decode_ENV_CTRL_2_86 = (decode_INSTRUCTION & 32'h00006014);
  assign _zz__zz_decode_ENV_CTRL_2_87 = 32'h00002010;
  assign _zz__zz_decode_ENV_CTRL_2_90 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_91) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_92 = {(_zz__zz_decode_ENV_CTRL_2_93 == _zz__zz_decode_ENV_CTRL_2_94),{_zz__zz_decode_ENV_CTRL_2_95,_zz__zz_decode_ENV_CTRL_2_96}};
  assign _zz__zz_decode_ENV_CTRL_2_98 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_99) == 32'h0);
  assign _zz__zz_decode_ENV_CTRL_2_100 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_102 = ({_zz__zz_decode_ENV_CTRL_2_103,{_zz__zz_decode_ENV_CTRL_2_104,_zz__zz_decode_ENV_CTRL_2_106}} != 3'b000);
  assign _zz__zz_decode_ENV_CTRL_2_108 = ({_zz__zz_decode_ENV_CTRL_2_109,_zz__zz_decode_ENV_CTRL_2_111} != 2'b00);
  assign _zz__zz_decode_ENV_CTRL_2_112 = {(_zz__zz_decode_ENV_CTRL_2_113 != _zz__zz_decode_ENV_CTRL_2_116),(_zz__zz_decode_ENV_CTRL_2_117 != _zz__zz_decode_ENV_CTRL_2_119)};
  assign _zz__zz_decode_ENV_CTRL_2_91 = 32'h00000044;
  assign _zz__zz_decode_ENV_CTRL_2_93 = (decode_INSTRUCTION & 32'h00000018);
  assign _zz__zz_decode_ENV_CTRL_2_94 = 32'h0;
  assign _zz__zz_decode_ENV_CTRL_2_95 = ((decode_INSTRUCTION & 32'h00006004) == 32'h00002000);
  assign _zz__zz_decode_ENV_CTRL_2_96 = ((decode_INSTRUCTION & 32'h00005004) == 32'h00001000);
  assign _zz__zz_decode_ENV_CTRL_2_99 = 32'h00000058;
  assign _zz__zz_decode_ENV_CTRL_2_103 = ((decode_INSTRUCTION & 32'h00000044) == 32'h00000040);
  assign _zz__zz_decode_ENV_CTRL_2_104 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_105) == 32'h00002010);
  assign _zz__zz_decode_ENV_CTRL_2_106 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_107) == 32'h40000030);
  assign _zz__zz_decode_ENV_CTRL_2_109 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_110) == 32'h00000004);
  assign _zz__zz_decode_ENV_CTRL_2_111 = _zz_decode_ENV_CTRL_3;
  assign _zz__zz_decode_ENV_CTRL_2_113 = {(_zz__zz_decode_ENV_CTRL_2_114 == _zz__zz_decode_ENV_CTRL_2_115),_zz_decode_ENV_CTRL_3};
  assign _zz__zz_decode_ENV_CTRL_2_116 = 2'b00;
  assign _zz__zz_decode_ENV_CTRL_2_117 = ((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2_118) == 32'h00001008);
  assign _zz__zz_decode_ENV_CTRL_2_119 = 1'b0;
  assign _zz__zz_decode_ENV_CTRL_2_105 = 32'h00002014;
  assign _zz__zz_decode_ENV_CTRL_2_107 = 32'h40004034;
  assign _zz__zz_decode_ENV_CTRL_2_110 = 32'h00000014;
  assign _zz__zz_decode_ENV_CTRL_2_114 = (decode_INSTRUCTION & 32'h00000044);
  assign _zz__zz_decode_ENV_CTRL_2_115 = 32'h00000004;
  assign _zz__zz_decode_ENV_CTRL_2_118 = 32'h00001048;
  always @(posedge clk) begin
    if(_zz_decode_RegFilePlugin_rs1Data) begin
      _zz_RegFilePlugin_regFile_port0 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress1];
    end
  end

  always @(posedge clk) begin
    if(_zz_decode_RegFilePlugin_rs2Data) begin
      _zz_RegFilePlugin_regFile_port1 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress2];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      RegFilePlugin_regFile[lastStageRegFileWrite_payload_address] <= lastStageRegFileWrite_payload_data;
    end
  end

  InstructionCache IBusCachedPlugin_cache (
    .io_flush                                 (IBusCachedPlugin_cache_io_flush                       ), //i
    .io_cpu_prefetch_isValid                  (IBusCachedPlugin_cache_io_cpu_prefetch_isValid        ), //i
    .io_cpu_prefetch_haltIt                   (IBusCachedPlugin_cache_io_cpu_prefetch_haltIt         ), //o
    .io_cpu_prefetch_pc                       (IBusCachedPlugin_iBusRsp_stages_0_input_payload       ), //i
    .io_cpu_fetch_isValid                     (IBusCachedPlugin_cache_io_cpu_fetch_isValid           ), //i
    .io_cpu_fetch_isStuck                     (IBusCachedPlugin_cache_io_cpu_fetch_isStuck           ), //i
    .io_cpu_fetch_isRemoved                   (IBusCachedPlugin_cache_io_cpu_fetch_isRemoved         ), //i
    .io_cpu_fetch_pc                          (IBusCachedPlugin_iBusRsp_stages_1_input_payload       ), //i
    .io_cpu_fetch_data                        (IBusCachedPlugin_cache_io_cpu_fetch_data              ), //o
    .io_cpu_fetch_mmuRsp_physicalAddress      (IBusCachedPlugin_mmuBus_rsp_physicalAddress           ), //i
    .io_cpu_fetch_mmuRsp_isIoAccess           (IBusCachedPlugin_mmuBus_rsp_isIoAccess                ), //i
    .io_cpu_fetch_mmuRsp_isPaging             (IBusCachedPlugin_mmuBus_rsp_isPaging                  ), //i
    .io_cpu_fetch_mmuRsp_allowRead            (IBusCachedPlugin_mmuBus_rsp_allowRead                 ), //i
    .io_cpu_fetch_mmuRsp_allowWrite           (IBusCachedPlugin_mmuBus_rsp_allowWrite                ), //i
    .io_cpu_fetch_mmuRsp_allowExecute         (IBusCachedPlugin_mmuBus_rsp_allowExecute              ), //i
    .io_cpu_fetch_mmuRsp_exception            (IBusCachedPlugin_mmuBus_rsp_exception                 ), //i
    .io_cpu_fetch_mmuRsp_refilling            (IBusCachedPlugin_mmuBus_rsp_refilling                 ), //i
    .io_cpu_fetch_mmuRsp_bypassTranslation    (IBusCachedPlugin_mmuBus_rsp_bypassTranslation         ), //i
    .io_cpu_fetch_physicalAddress             (IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress   ), //o
    .io_cpu_decode_isValid                    (IBusCachedPlugin_cache_io_cpu_decode_isValid          ), //i
    .io_cpu_decode_isStuck                    (IBusCachedPlugin_cache_io_cpu_decode_isStuck          ), //i
    .io_cpu_decode_pc                         (IBusCachedPlugin_iBusRsp_stages_2_input_payload       ), //i
    .io_cpu_decode_physicalAddress            (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress  ), //o
    .io_cpu_decode_data                       (IBusCachedPlugin_cache_io_cpu_decode_data             ), //o
    .io_cpu_decode_cacheMiss                  (IBusCachedPlugin_cache_io_cpu_decode_cacheMiss        ), //o
    .io_cpu_decode_error                      (IBusCachedPlugin_cache_io_cpu_decode_error            ), //o
    .io_cpu_decode_mmuRefilling               (IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling     ), //o
    .io_cpu_decode_mmuException               (IBusCachedPlugin_cache_io_cpu_decode_mmuException     ), //o
    .io_cpu_decode_isUser                     (IBusCachedPlugin_cache_io_cpu_decode_isUser           ), //i
    .io_cpu_fill_valid                        (IBusCachedPlugin_cache_io_cpu_fill_valid              ), //i
    .io_cpu_fill_payload                      (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress  ), //i
    .io_mem_cmd_valid                         (IBusCachedPlugin_cache_io_mem_cmd_valid               ), //o
    .io_mem_cmd_ready                         (iBus_cmd_ready                                        ), //i
    .io_mem_cmd_payload_address               (IBusCachedPlugin_cache_io_mem_cmd_payload_address     ), //o
    .io_mem_cmd_payload_size                  (IBusCachedPlugin_cache_io_mem_cmd_payload_size        ), //o
    .io_mem_rsp_valid                         (iBus_rsp_valid                                        ), //i
    .io_mem_rsp_payload_data                  (iBus_rsp_payload_data                                 ), //i
    .io_mem_rsp_payload_error                 (iBus_rsp_payload_error                                ), //i
    ._zz_when_Fetcher_l398                    (switch_Fetcher_l362                                   ), //i
    ._zz_io_cpu_fetch_data_regNextWhen        (IBusCachedPlugin_injectionPort_payload                ), //i
    .clk                                      (clk                                                   ), //i
    .reset                                    (reset                                                 )  //i
  );
  
  always @(*) begin
    case(_zz_memory_to_writeBack_ENV_CTRL)
      2'b00 : _zz_memory_to_writeBack_ENV_CTRL_string = "NONE ";
      2'b01 : _zz_memory_to_writeBack_ENV_CTRL_string = "XRET ";
      2'b10 : _zz_memory_to_writeBack_ENV_CTRL_string = "ECALL";
      default : _zz_memory_to_writeBack_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_ENV_CTRL_1)
      2'b00 : _zz_memory_to_writeBack_ENV_CTRL_1_string = "NONE ";
      2'b01 : _zz_memory_to_writeBack_ENV_CTRL_1_string = "XRET ";
      2'b10 : _zz_memory_to_writeBack_ENV_CTRL_1_string = "ECALL";
      default : _zz_memory_to_writeBack_ENV_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_ENV_CTRL)
      2'b00 : _zz_execute_to_memory_ENV_CTRL_string = "NONE ";
      2'b01 : _zz_execute_to_memory_ENV_CTRL_string = "XRET ";
      2'b10 : _zz_execute_to_memory_ENV_CTRL_string = "ECALL";
      default : _zz_execute_to_memory_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_ENV_CTRL_1)
      2'b00 : _zz_execute_to_memory_ENV_CTRL_1_string = "NONE ";
      2'b01 : _zz_execute_to_memory_ENV_CTRL_1_string = "XRET ";
      2'b10 : _zz_execute_to_memory_ENV_CTRL_1_string = "ECALL";
      default : _zz_execute_to_memory_ENV_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_ENV_CTRL)
      2'b00 : decode_ENV_CTRL_string = "NONE ";
      2'b01 : decode_ENV_CTRL_string = "XRET ";
      2'b10 : decode_ENV_CTRL_string = "ECALL";
      default : decode_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL)
      2'b00 : _zz_decode_ENV_CTRL_string = "NONE ";
      2'b01 : _zz_decode_ENV_CTRL_string = "XRET ";
      2'b10 : _zz_decode_ENV_CTRL_string = "ECALL";
      default : _zz_decode_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ENV_CTRL)
      2'b00 : _zz_decode_to_execute_ENV_CTRL_string = "NONE ";
      2'b01 : _zz_decode_to_execute_ENV_CTRL_string = "XRET ";
      2'b10 : _zz_decode_to_execute_ENV_CTRL_string = "ECALL";
      default : _zz_decode_to_execute_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ENV_CTRL_1)
      2'b00 : _zz_decode_to_execute_ENV_CTRL_1_string = "NONE ";
      2'b01 : _zz_decode_to_execute_ENV_CTRL_1_string = "XRET ";
      2'b10 : _zz_decode_to_execute_ENV_CTRL_1_string = "ECALL";
      default : _zz_decode_to_execute_ENV_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_BRANCH_CTRL)
      2'b00 : decode_BRANCH_CTRL_string = "INC ";
      2'b01 : decode_BRANCH_CTRL_string = "B   ";
      2'b10 : decode_BRANCH_CTRL_string = "JAL ";
      2'b11 : decode_BRANCH_CTRL_string = "JALR";
      default : decode_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL)
      2'b00 : _zz_decode_BRANCH_CTRL_string = "INC ";
      2'b01 : _zz_decode_BRANCH_CTRL_string = "B   ";
      2'b10 : _zz_decode_BRANCH_CTRL_string = "JAL ";
      2'b11 : _zz_decode_BRANCH_CTRL_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_BRANCH_CTRL)
      2'b00 : _zz_decode_to_execute_BRANCH_CTRL_string = "INC ";
      2'b01 : _zz_decode_to_execute_BRANCH_CTRL_string = "B   ";
      2'b10 : _zz_decode_to_execute_BRANCH_CTRL_string = "JAL ";
      2'b11 : _zz_decode_to_execute_BRANCH_CTRL_string = "JALR";
      default : _zz_decode_to_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_BRANCH_CTRL_1)
      2'b00 : _zz_decode_to_execute_BRANCH_CTRL_1_string = "INC ";
      2'b01 : _zz_decode_to_execute_BRANCH_CTRL_1_string = "B   ";
      2'b10 : _zz_decode_to_execute_BRANCH_CTRL_1_string = "JAL ";
      2'b11 : _zz_decode_to_execute_BRANCH_CTRL_1_string = "JALR";
      default : _zz_decode_to_execute_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(decode_SHIFT_CTRL)
      2'b00 : decode_SHIFT_CTRL_string = "DISABLE_1";
      2'b01 : decode_SHIFT_CTRL_string = "SLL_1    ";
      2'b10 : decode_SHIFT_CTRL_string = "SRL_1    ";
      2'b11 : decode_SHIFT_CTRL_string = "SRA_1    ";
      default : decode_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL)
      2'b00 : _zz_decode_SHIFT_CTRL_string = "DISABLE_1";
      2'b01 : _zz_decode_SHIFT_CTRL_string = "SLL_1    ";
      2'b10 : _zz_decode_SHIFT_CTRL_string = "SRL_1    ";
      2'b11 : _zz_decode_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SHIFT_CTRL)
      2'b00 : _zz_decode_to_execute_SHIFT_CTRL_string = "DISABLE_1";
      2'b01 : _zz_decode_to_execute_SHIFT_CTRL_string = "SLL_1    ";
      2'b10 : _zz_decode_to_execute_SHIFT_CTRL_string = "SRL_1    ";
      2'b11 : _zz_decode_to_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_decode_to_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SHIFT_CTRL_1)
      2'b00 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "DISABLE_1";
      2'b01 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SLL_1    ";
      2'b10 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SRL_1    ";
      2'b11 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_decode_to_execute_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_ALU_BITWISE_CTRL)
      2'b00 : decode_ALU_BITWISE_CTRL_string = "XOR_1";
      2'b01 : decode_ALU_BITWISE_CTRL_string = "OR_1 ";
      2'b10 : decode_ALU_BITWISE_CTRL_string = "AND_1";
      default : decode_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL)
      2'b00 : _zz_decode_ALU_BITWISE_CTRL_string = "XOR_1";
      2'b01 : _zz_decode_ALU_BITWISE_CTRL_string = "OR_1 ";
      2'b10 : _zz_decode_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_BITWISE_CTRL)
      2'b00 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      2'b01 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      2'b10 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_BITWISE_CTRL_1)
      2'b00 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "XOR_1";
      2'b01 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      2'b10 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_SRC2_CTRL)
      2'b00 : decode_SRC2_CTRL_string = "RS ";
      2'b01 : decode_SRC2_CTRL_string = "IMI";
      2'b10 : decode_SRC2_CTRL_string = "IMS";
      2'b11 : decode_SRC2_CTRL_string = "PC ";
      default : decode_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL)
      2'b00 : _zz_decode_SRC2_CTRL_string = "RS ";
      2'b01 : _zz_decode_SRC2_CTRL_string = "IMI";
      2'b10 : _zz_decode_SRC2_CTRL_string = "IMS";
      2'b11 : _zz_decode_SRC2_CTRL_string = "PC ";
      default : _zz_decode_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SRC2_CTRL)
      2'b00 : _zz_decode_to_execute_SRC2_CTRL_string = "RS ";
      2'b01 : _zz_decode_to_execute_SRC2_CTRL_string = "IMI";
      2'b10 : _zz_decode_to_execute_SRC2_CTRL_string = "IMS";
      2'b11 : _zz_decode_to_execute_SRC2_CTRL_string = "PC ";
      default : _zz_decode_to_execute_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SRC2_CTRL_1)
      2'b00 : _zz_decode_to_execute_SRC2_CTRL_1_string = "RS ";
      2'b01 : _zz_decode_to_execute_SRC2_CTRL_1_string = "IMI";
      2'b10 : _zz_decode_to_execute_SRC2_CTRL_1_string = "IMS";
      2'b11 : _zz_decode_to_execute_SRC2_CTRL_1_string = "PC ";
      default : _zz_decode_to_execute_SRC2_CTRL_1_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_ALU_CTRL)
      2'b00 : decode_ALU_CTRL_string = "ADD_SUB ";
      2'b01 : decode_ALU_CTRL_string = "SLT_SLTU";
      2'b10 : decode_ALU_CTRL_string = "BITWISE ";
      default : decode_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL)
      2'b00 : _zz_decode_ALU_CTRL_string = "ADD_SUB ";
      2'b01 : _zz_decode_ALU_CTRL_string = "SLT_SLTU";
      2'b10 : _zz_decode_ALU_CTRL_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_CTRL)
      2'b00 : _zz_decode_to_execute_ALU_CTRL_string = "ADD_SUB ";
      2'b01 : _zz_decode_to_execute_ALU_CTRL_string = "SLT_SLTU";
      2'b10 : _zz_decode_to_execute_ALU_CTRL_string = "BITWISE ";
      default : _zz_decode_to_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_CTRL_1)
      2'b00 : _zz_decode_to_execute_ALU_CTRL_1_string = "ADD_SUB ";
      2'b01 : _zz_decode_to_execute_ALU_CTRL_1_string = "SLT_SLTU";
      2'b10 : _zz_decode_to_execute_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_decode_to_execute_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_SRC1_CTRL)
      2'b00 : decode_SRC1_CTRL_string = "RS          ";
      2'b01 : decode_SRC1_CTRL_string = "IMU         ";
      2'b10 : decode_SRC1_CTRL_string = "PC_INCREMENT";
      2'b11 : decode_SRC1_CTRL_string = "URS1        ";
      default : decode_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL)
      2'b00 : _zz_decode_SRC1_CTRL_string = "RS          ";
      2'b01 : _zz_decode_SRC1_CTRL_string = "IMU         ";
      2'b10 : _zz_decode_SRC1_CTRL_string = "PC_INCREMENT";
      2'b11 : _zz_decode_SRC1_CTRL_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SRC1_CTRL)
      2'b00 : _zz_decode_to_execute_SRC1_CTRL_string = "RS          ";
      2'b01 : _zz_decode_to_execute_SRC1_CTRL_string = "IMU         ";
      2'b10 : _zz_decode_to_execute_SRC1_CTRL_string = "PC_INCREMENT";
      2'b11 : _zz_decode_to_execute_SRC1_CTRL_string = "URS1        ";
      default : _zz_decode_to_execute_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SRC1_CTRL_1)
      2'b00 : _zz_decode_to_execute_SRC1_CTRL_1_string = "RS          ";
      2'b01 : _zz_decode_to_execute_SRC1_CTRL_1_string = "IMU         ";
      2'b10 : _zz_decode_to_execute_SRC1_CTRL_1_string = "PC_INCREMENT";
      2'b11 : _zz_decode_to_execute_SRC1_CTRL_1_string = "URS1        ";
      default : _zz_decode_to_execute_SRC1_CTRL_1_string = "????????????";
    endcase
  end
  always @(*) begin
    case(memory_ENV_CTRL)
      2'b00 : memory_ENV_CTRL_string = "NONE ";
      2'b01 : memory_ENV_CTRL_string = "XRET ";
      2'b10 : memory_ENV_CTRL_string = "ECALL";
      default : memory_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_ENV_CTRL)
      2'b00 : _zz_memory_ENV_CTRL_string = "NONE ";
      2'b01 : _zz_memory_ENV_CTRL_string = "XRET ";
      2'b10 : _zz_memory_ENV_CTRL_string = "ECALL";
      default : _zz_memory_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ENV_CTRL)
      2'b00 : execute_ENV_CTRL_string = "NONE ";
      2'b01 : execute_ENV_CTRL_string = "XRET ";
      2'b10 : execute_ENV_CTRL_string = "ECALL";
      default : execute_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ENV_CTRL)
      2'b00 : _zz_execute_ENV_CTRL_string = "NONE ";
      2'b01 : _zz_execute_ENV_CTRL_string = "XRET ";
      2'b10 : _zz_execute_ENV_CTRL_string = "ECALL";
      default : _zz_execute_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(writeBack_ENV_CTRL)
      2'b00 : writeBack_ENV_CTRL_string = "NONE ";
      2'b01 : writeBack_ENV_CTRL_string = "XRET ";
      2'b10 : writeBack_ENV_CTRL_string = "ECALL";
      default : writeBack_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_writeBack_ENV_CTRL)
      2'b00 : _zz_writeBack_ENV_CTRL_string = "NONE ";
      2'b01 : _zz_writeBack_ENV_CTRL_string = "XRET ";
      2'b10 : _zz_writeBack_ENV_CTRL_string = "ECALL";
      default : _zz_writeBack_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_BRANCH_CTRL)
      2'b00 : execute_BRANCH_CTRL_string = "INC ";
      2'b01 : execute_BRANCH_CTRL_string = "B   ";
      2'b10 : execute_BRANCH_CTRL_string = "JAL ";
      2'b11 : execute_BRANCH_CTRL_string = "JALR";
      default : execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_BRANCH_CTRL)
      2'b00 : _zz_execute_BRANCH_CTRL_string = "INC ";
      2'b01 : _zz_execute_BRANCH_CTRL_string = "B   ";
      2'b10 : _zz_execute_BRANCH_CTRL_string = "JAL ";
      2'b11 : _zz_execute_BRANCH_CTRL_string = "JALR";
      default : _zz_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_SHIFT_CTRL)
      2'b00 : execute_SHIFT_CTRL_string = "DISABLE_1";
      2'b01 : execute_SHIFT_CTRL_string = "SLL_1    ";
      2'b10 : execute_SHIFT_CTRL_string = "SRL_1    ";
      2'b11 : execute_SHIFT_CTRL_string = "SRA_1    ";
      default : execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_SHIFT_CTRL)
      2'b00 : _zz_execute_SHIFT_CTRL_string = "DISABLE_1";
      2'b01 : _zz_execute_SHIFT_CTRL_string = "SLL_1    ";
      2'b10 : _zz_execute_SHIFT_CTRL_string = "SRL_1    ";
      2'b11 : _zz_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_SRC2_CTRL)
      2'b00 : execute_SRC2_CTRL_string = "RS ";
      2'b01 : execute_SRC2_CTRL_string = "IMI";
      2'b10 : execute_SRC2_CTRL_string = "IMS";
      2'b11 : execute_SRC2_CTRL_string = "PC ";
      default : execute_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_execute_SRC2_CTRL)
      2'b00 : _zz_execute_SRC2_CTRL_string = "RS ";
      2'b01 : _zz_execute_SRC2_CTRL_string = "IMI";
      2'b10 : _zz_execute_SRC2_CTRL_string = "IMS";
      2'b11 : _zz_execute_SRC2_CTRL_string = "PC ";
      default : _zz_execute_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_SRC1_CTRL)
      2'b00 : execute_SRC1_CTRL_string = "RS          ";
      2'b01 : execute_SRC1_CTRL_string = "IMU         ";
      2'b10 : execute_SRC1_CTRL_string = "PC_INCREMENT";
      2'b11 : execute_SRC1_CTRL_string = "URS1        ";
      default : execute_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_SRC1_CTRL)
      2'b00 : _zz_execute_SRC1_CTRL_string = "RS          ";
      2'b01 : _zz_execute_SRC1_CTRL_string = "IMU         ";
      2'b10 : _zz_execute_SRC1_CTRL_string = "PC_INCREMENT";
      2'b11 : _zz_execute_SRC1_CTRL_string = "URS1        ";
      default : _zz_execute_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(execute_ALU_CTRL)
      2'b00 : execute_ALU_CTRL_string = "ADD_SUB ";
      2'b01 : execute_ALU_CTRL_string = "SLT_SLTU";
      2'b10 : execute_ALU_CTRL_string = "BITWISE ";
      default : execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ALU_CTRL)
      2'b00 : _zz_execute_ALU_CTRL_string = "ADD_SUB ";
      2'b01 : _zz_execute_ALU_CTRL_string = "SLT_SLTU";
      2'b10 : _zz_execute_ALU_CTRL_string = "BITWISE ";
      default : _zz_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_ALU_BITWISE_CTRL)
      2'b00 : execute_ALU_BITWISE_CTRL_string = "XOR_1";
      2'b01 : execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      2'b10 : execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ALU_BITWISE_CTRL)
      2'b00 : _zz_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      2'b01 : _zz_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      2'b10 : _zz_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL_1)
      2'b00 : _zz_decode_ENV_CTRL_1_string = "NONE ";
      2'b01 : _zz_decode_ENV_CTRL_1_string = "XRET ";
      2'b10 : _zz_decode_ENV_CTRL_1_string = "ECALL";
      default : _zz_decode_ENV_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL_1)
      2'b00 : _zz_decode_BRANCH_CTRL_1_string = "INC ";
      2'b01 : _zz_decode_BRANCH_CTRL_1_string = "B   ";
      2'b10 : _zz_decode_BRANCH_CTRL_1_string = "JAL ";
      2'b11 : _zz_decode_BRANCH_CTRL_1_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL_1)
      2'b00 : _zz_decode_SHIFT_CTRL_1_string = "DISABLE_1";
      2'b01 : _zz_decode_SHIFT_CTRL_1_string = "SLL_1    ";
      2'b10 : _zz_decode_SHIFT_CTRL_1_string = "SRL_1    ";
      2'b11 : _zz_decode_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL_1)
      2'b00 : _zz_decode_ALU_BITWISE_CTRL_1_string = "XOR_1";
      2'b01 : _zz_decode_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      2'b10 : _zz_decode_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL_1)
      2'b00 : _zz_decode_SRC2_CTRL_1_string = "RS ";
      2'b01 : _zz_decode_SRC2_CTRL_1_string = "IMI";
      2'b10 : _zz_decode_SRC2_CTRL_1_string = "IMS";
      2'b11 : _zz_decode_SRC2_CTRL_1_string = "PC ";
      default : _zz_decode_SRC2_CTRL_1_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL_1)
      2'b00 : _zz_decode_ALU_CTRL_1_string = "ADD_SUB ";
      2'b01 : _zz_decode_ALU_CTRL_1_string = "SLT_SLTU";
      2'b10 : _zz_decode_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL_1)
      2'b00 : _zz_decode_SRC1_CTRL_1_string = "RS          ";
      2'b01 : _zz_decode_SRC1_CTRL_1_string = "IMU         ";
      2'b10 : _zz_decode_SRC1_CTRL_1_string = "PC_INCREMENT";
      2'b11 : _zz_decode_SRC1_CTRL_1_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_1_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL_2)
      2'b00 : _zz_decode_SRC1_CTRL_2_string = "RS          ";
      2'b01 : _zz_decode_SRC1_CTRL_2_string = "IMU         ";
      2'b10 : _zz_decode_SRC1_CTRL_2_string = "PC_INCREMENT";
      2'b11 : _zz_decode_SRC1_CTRL_2_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_2_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL_2)
      2'b00 : _zz_decode_ALU_CTRL_2_string = "ADD_SUB ";
      2'b01 : _zz_decode_ALU_CTRL_2_string = "SLT_SLTU";
      2'b10 : _zz_decode_ALU_CTRL_2_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL_2)
      2'b00 : _zz_decode_SRC2_CTRL_2_string = "RS ";
      2'b01 : _zz_decode_SRC2_CTRL_2_string = "IMI";
      2'b10 : _zz_decode_SRC2_CTRL_2_string = "IMS";
      2'b11 : _zz_decode_SRC2_CTRL_2_string = "PC ";
      default : _zz_decode_SRC2_CTRL_2_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL_2)
      2'b00 : _zz_decode_ALU_BITWISE_CTRL_2_string = "XOR_1";
      2'b01 : _zz_decode_ALU_BITWISE_CTRL_2_string = "OR_1 ";
      2'b10 : _zz_decode_ALU_BITWISE_CTRL_2_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL_2)
      2'b00 : _zz_decode_SHIFT_CTRL_2_string = "DISABLE_1";
      2'b01 : _zz_decode_SHIFT_CTRL_2_string = "SLL_1    ";
      2'b10 : _zz_decode_SHIFT_CTRL_2_string = "SRL_1    ";
      2'b11 : _zz_decode_SHIFT_CTRL_2_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_2_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL_2)
      2'b00 : _zz_decode_BRANCH_CTRL_2_string = "INC ";
      2'b01 : _zz_decode_BRANCH_CTRL_2_string = "B   ";
      2'b10 : _zz_decode_BRANCH_CTRL_2_string = "JAL ";
      2'b11 : _zz_decode_BRANCH_CTRL_2_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL_7)
      2'b00 : _zz_decode_ENV_CTRL_7_string = "NONE ";
      2'b01 : _zz_decode_ENV_CTRL_7_string = "XRET ";
      2'b10 : _zz_decode_ENV_CTRL_7_string = "ECALL";
      default : _zz_decode_ENV_CTRL_7_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_SRC1_CTRL)
      2'b00 : decode_to_execute_SRC1_CTRL_string = "RS          ";
      2'b01 : decode_to_execute_SRC1_CTRL_string = "IMU         ";
      2'b10 : decode_to_execute_SRC1_CTRL_string = "PC_INCREMENT";
      2'b11 : decode_to_execute_SRC1_CTRL_string = "URS1        ";
      default : decode_to_execute_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ALU_CTRL)
      2'b00 : decode_to_execute_ALU_CTRL_string = "ADD_SUB ";
      2'b01 : decode_to_execute_ALU_CTRL_string = "SLT_SLTU";
      2'b10 : decode_to_execute_ALU_CTRL_string = "BITWISE ";
      default : decode_to_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_SRC2_CTRL)
      2'b00 : decode_to_execute_SRC2_CTRL_string = "RS ";
      2'b01 : decode_to_execute_SRC2_CTRL_string = "IMI";
      2'b10 : decode_to_execute_SRC2_CTRL_string = "IMS";
      2'b11 : decode_to_execute_SRC2_CTRL_string = "PC ";
      default : decode_to_execute_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ALU_BITWISE_CTRL)
      2'b00 : decode_to_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      2'b01 : decode_to_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      2'b10 : decode_to_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : decode_to_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_SHIFT_CTRL)
      2'b00 : decode_to_execute_SHIFT_CTRL_string = "DISABLE_1";
      2'b01 : decode_to_execute_SHIFT_CTRL_string = "SLL_1    ";
      2'b10 : decode_to_execute_SHIFT_CTRL_string = "SRL_1    ";
      2'b11 : decode_to_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : decode_to_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_BRANCH_CTRL)
      2'b00 : decode_to_execute_BRANCH_CTRL_string = "INC ";
      2'b01 : decode_to_execute_BRANCH_CTRL_string = "B   ";
      2'b10 : decode_to_execute_BRANCH_CTRL_string = "JAL ";
      2'b11 : decode_to_execute_BRANCH_CTRL_string = "JALR";
      default : decode_to_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ENV_CTRL)
      2'b00 : decode_to_execute_ENV_CTRL_string = "NONE ";
      2'b01 : decode_to_execute_ENV_CTRL_string = "XRET ";
      2'b10 : decode_to_execute_ENV_CTRL_string = "ECALL";
      default : decode_to_execute_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_ENV_CTRL)
      2'b00 : execute_to_memory_ENV_CTRL_string = "NONE ";
      2'b01 : execute_to_memory_ENV_CTRL_string = "XRET ";
      2'b10 : execute_to_memory_ENV_CTRL_string = "ECALL";
      default : execute_to_memory_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(memory_to_writeBack_ENV_CTRL)
      2'b00 : memory_to_writeBack_ENV_CTRL_string = "NONE ";
      2'b01 : memory_to_writeBack_ENV_CTRL_string = "XRET ";
      2'b10 : memory_to_writeBack_ENV_CTRL_string = "ECALL";
      default : memory_to_writeBack_ENV_CTRL_string = "?????";
    endcase
  end
  

  assign memory_MEMORY_READ_DATA = dBus_rsp_data;
  assign execute_BRANCH_CALC = {execute_BranchPlugin_branchAdder[31 : 1],1'b0};
  assign execute_BRANCH_DO = _zz_execute_BRANCH_DO_1;
  assign writeBack_REGFILE_WRITE_DATA = memory_to_writeBack_REGFILE_WRITE_DATA;
  assign execute_REGFILE_WRITE_DATA = _zz_execute_REGFILE_WRITE_DATA;
  assign memory_MEMORY_ADDRESS_LOW = execute_to_memory_MEMORY_ADDRESS_LOW;
  assign execute_MEMORY_ADDRESS_LOW = dBus_cmd_payload_address[1 : 0];
  assign decode_DO_EBREAK = (((! DebugPlugin_haltIt) && (decode_IS_EBREAK || 1'b0)) && DebugPlugin_allowEBreak);
  assign decode_CSR_READ_OPCODE = (decode_INSTRUCTION[13 : 7] != 7'h20);
  assign decode_CSR_WRITE_OPCODE = (! (((decode_INSTRUCTION[14 : 13] == 2'b01) && (decode_INSTRUCTION[19 : 15] == 5'h0)) || ((decode_INSTRUCTION[14 : 13] == 2'b11) && (decode_INSTRUCTION[19 : 15] == 5'h0))));
  assign decode_SRC2_FORCE_ZERO = (decode_SRC_ADD_ZERO && (! decode_SRC_USE_SUB_LESS));
  assign decode_RS2 = decode_RegFilePlugin_rs2Data;
  assign decode_RS1 = decode_RegFilePlugin_rs1Data;
  assign _zz_memory_to_writeBack_ENV_CTRL = _zz_memory_to_writeBack_ENV_CTRL_1;
  assign _zz_execute_to_memory_ENV_CTRL = _zz_execute_to_memory_ENV_CTRL_1;
  assign decode_ENV_CTRL = _zz_decode_ENV_CTRL;
  assign _zz_decode_to_execute_ENV_CTRL = _zz_decode_to_execute_ENV_CTRL_1;
  assign decode_IS_CSR = _zz_decode_ENV_CTRL_2[24];
  assign decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL = _zz_decode_to_execute_BRANCH_CTRL_1;
  assign decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL = _zz_decode_to_execute_SHIFT_CTRL_1;
  assign decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL = _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  assign decode_SRC_LESS_UNSIGNED = _zz_decode_ENV_CTRL_2[16];
  assign decode_MEMORY_STORE = _zz_decode_ENV_CTRL_2[13];
  assign execute_BYPASSABLE_MEMORY_STAGE = decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  assign decode_BYPASSABLE_MEMORY_STAGE = _zz_decode_ENV_CTRL_2[12];
  assign decode_BYPASSABLE_EXECUTE_STAGE = _zz_decode_ENV_CTRL_2[11];
  assign decode_SRC2_CTRL = _zz_decode_SRC2_CTRL;
  assign _zz_decode_to_execute_SRC2_CTRL = _zz_decode_to_execute_SRC2_CTRL_1;
  assign decode_ALU_CTRL = _zz_decode_ALU_CTRL;
  assign _zz_decode_to_execute_ALU_CTRL = _zz_decode_to_execute_ALU_CTRL_1;
  assign decode_MEMORY_ENABLE = _zz_decode_ENV_CTRL_2[4];
  assign decode_SRC1_CTRL = _zz_decode_SRC1_CTRL;
  assign _zz_decode_to_execute_SRC1_CTRL = _zz_decode_to_execute_SRC1_CTRL_1;
  assign writeBack_FORMAL_PC_NEXT = memory_to_writeBack_FORMAL_PC_NEXT;
  assign memory_FORMAL_PC_NEXT = execute_to_memory_FORMAL_PC_NEXT;
  assign execute_FORMAL_PC_NEXT = decode_to_execute_FORMAL_PC_NEXT;
  assign decode_FORMAL_PC_NEXT = (decode_PC + 32'h00000004);
  assign memory_PC = execute_to_memory_PC;
  assign execute_DO_EBREAK = decode_to_execute_DO_EBREAK;
  assign decode_IS_EBREAK = _zz_decode_ENV_CTRL_2[27];
  assign execute_CSR_READ_OPCODE = decode_to_execute_CSR_READ_OPCODE;
  assign execute_CSR_WRITE_OPCODE = decode_to_execute_CSR_WRITE_OPCODE;
  assign execute_IS_CSR = decode_to_execute_IS_CSR;
  assign memory_ENV_CTRL = _zz_memory_ENV_CTRL;
  assign execute_ENV_CTRL = _zz_execute_ENV_CTRL;
  assign writeBack_ENV_CTRL = _zz_writeBack_ENV_CTRL;
  assign memory_BRANCH_CALC = execute_to_memory_BRANCH_CALC;
  assign memory_BRANCH_DO = execute_to_memory_BRANCH_DO;
  assign execute_PC = decode_to_execute_PC;
  assign execute_RS1 = decode_to_execute_RS1;
  assign execute_BRANCH_CTRL = _zz_execute_BRANCH_CTRL;
  assign decode_RS2_USE = _zz_decode_ENV_CTRL_2[15];
  assign decode_RS1_USE = _zz_decode_ENV_CTRL_2[5];
  assign execute_REGFILE_WRITE_VALID = decode_to_execute_REGFILE_WRITE_VALID;
  assign execute_BYPASSABLE_EXECUTE_STAGE = decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  assign memory_REGFILE_WRITE_VALID = execute_to_memory_REGFILE_WRITE_VALID;
  assign memory_INSTRUCTION = execute_to_memory_INSTRUCTION;
  assign memory_BYPASSABLE_MEMORY_STAGE = execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  assign writeBack_REGFILE_WRITE_VALID = memory_to_writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    _zz_execute_to_memory_REGFILE_WRITE_DATA = execute_REGFILE_WRITE_DATA;
    if(when_ShiftPlugins_l169) begin
      _zz_execute_to_memory_REGFILE_WRITE_DATA = _zz_execute_to_memory_REGFILE_WRITE_DATA_1;
    end
    if(when_CsrPlugin_l1176) begin
      _zz_execute_to_memory_REGFILE_WRITE_DATA = CsrPlugin_csrMapping_readDataSignal;
    end
  end

  assign execute_SHIFT_CTRL = _zz_execute_SHIFT_CTRL;
  assign execute_SRC_LESS_UNSIGNED = decode_to_execute_SRC_LESS_UNSIGNED;
  assign execute_SRC2_FORCE_ZERO = decode_to_execute_SRC2_FORCE_ZERO;
  assign execute_SRC_USE_SUB_LESS = decode_to_execute_SRC_USE_SUB_LESS;
  assign _zz_execute_SRC2 = execute_PC;
  assign execute_SRC2_CTRL = _zz_execute_SRC2_CTRL;
  assign execute_SRC1_CTRL = _zz_execute_SRC1_CTRL;
  assign decode_SRC_USE_SUB_LESS = _zz_decode_ENV_CTRL_2[3];
  assign decode_SRC_ADD_ZERO = _zz_decode_ENV_CTRL_2[19];
  assign execute_SRC_ADD_SUB = execute_SrcPlugin_addSub;
  assign execute_SRC_LESS = execute_SrcPlugin_less;
  assign execute_ALU_CTRL = _zz_execute_ALU_CTRL;
  assign execute_SRC2 = _zz_execute_SRC2_5;
  assign execute_SRC1 = _zz_execute_SRC1;
  assign execute_ALU_BITWISE_CTRL = _zz_execute_ALU_BITWISE_CTRL;
  assign _zz_lastStageRegFileWrite_payload_address = writeBack_INSTRUCTION;
  assign _zz_lastStageRegFileWrite_valid = writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    _zz_1 = 1'b0;
    if(lastStageRegFileWrite_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign decode_INSTRUCTION_ANTICIPATED = (decode_arbitration_isStuck ? decode_INSTRUCTION : IBusCachedPlugin_cache_io_cpu_fetch_data);
  always @(*) begin
    decode_REGFILE_WRITE_VALID = _zz_decode_ENV_CTRL_2[10];
    if(when_RegFilePlugin_l63) begin
      decode_REGFILE_WRITE_VALID = 1'b0;
    end
  end

  assign decode_LEGAL_INSTRUCTION = ({((decode_INSTRUCTION & 32'h0000005f) == 32'h00000017),{((decode_INSTRUCTION & 32'h0000007f) == 32'h0000006f),{((decode_INSTRUCTION & 32'h0000106f) == 32'h00000003),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION) == 32'h00001073),{(_zz_decode_LEGAL_INSTRUCTION_1 == _zz_decode_LEGAL_INSTRUCTION_2),{_zz_decode_LEGAL_INSTRUCTION_3,{_zz_decode_LEGAL_INSTRUCTION_4,_zz_decode_LEGAL_INSTRUCTION_5}}}}}}} != 20'h0);
  assign writeBack_MEMORY_STORE = memory_to_writeBack_MEMORY_STORE;
  always @(*) begin
    _zz_lastStageRegFileWrite_payload_data = writeBack_REGFILE_WRITE_DATA;
    if(when_DBusSimplePlugin_l558) begin
      _zz_lastStageRegFileWrite_payload_data = writeBack_DBusSimplePlugin_rspFormated;
    end
  end

  assign writeBack_MEMORY_ENABLE = memory_to_writeBack_MEMORY_ENABLE;
  assign writeBack_MEMORY_ADDRESS_LOW = memory_to_writeBack_MEMORY_ADDRESS_LOW;
  assign writeBack_MEMORY_READ_DATA = memory_to_writeBack_MEMORY_READ_DATA;
  assign memory_ALIGNEMENT_FAULT = execute_to_memory_ALIGNEMENT_FAULT;
  assign memory_REGFILE_WRITE_DATA = execute_to_memory_REGFILE_WRITE_DATA;
  assign memory_MEMORY_STORE = execute_to_memory_MEMORY_STORE;
  assign memory_MEMORY_ENABLE = execute_to_memory_MEMORY_ENABLE;
  assign execute_SRC_ADD = execute_SrcPlugin_addSub;
  assign execute_RS2 = decode_to_execute_RS2;
  assign execute_INSTRUCTION = decode_to_execute_INSTRUCTION;
  assign execute_MEMORY_STORE = decode_to_execute_MEMORY_STORE;
  assign execute_MEMORY_ENABLE = decode_to_execute_MEMORY_ENABLE;
  assign execute_ALIGNEMENT_FAULT = (((dBus_cmd_payload_size == 2'b10) && (dBus_cmd_payload_address[1 : 0] != 2'b00)) || ((dBus_cmd_payload_size == 2'b01) && (dBus_cmd_payload_address[0 : 0] != 1'b0)));
  assign decode_FLUSH_ALL = _zz_decode_ENV_CTRL_2[0];
  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_4 = IBusCachedPlugin_rsp_issueDetected_3;
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_rsp_issueDetected_4 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_3 = IBusCachedPlugin_rsp_issueDetected_2;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_rsp_issueDetected_3 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_2 = IBusCachedPlugin_rsp_issueDetected_1;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_rsp_issueDetected_2 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_1 = IBusCachedPlugin_rsp_issueDetected;
    if(when_IBusCachedPlugin_l239) begin
      IBusCachedPlugin_rsp_issueDetected_1 = 1'b1;
    end
  end

  assign decode_INSTRUCTION = IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  always @(*) begin
    _zz_memory_to_writeBack_FORMAL_PC_NEXT = memory_FORMAL_PC_NEXT;
    if(BranchPlugin_jumpInterface_valid) begin
      _zz_memory_to_writeBack_FORMAL_PC_NEXT = BranchPlugin_jumpInterface_payload;
    end
  end

  assign decode_PC = IBusCachedPlugin_iBusRsp_output_payload_pc;
  assign writeBack_PC = memory_to_writeBack_PC;
  assign writeBack_INSTRUCTION = memory_to_writeBack_INSTRUCTION;
  always @(*) begin
    decode_arbitration_haltItself = 1'b0;
    case(switch_Fetcher_l362)
      3'b010 : begin
        decode_arbitration_haltItself = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    decode_arbitration_haltByOther = 1'b0;
    if(when_HazardSimplePlugin_l113) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    if(CsrPlugin_pipelineLiberator_active) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    if(when_CsrPlugin_l1116) begin
      decode_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    decode_arbitration_removeIt = 1'b0;
    if(_zz_when) begin
      decode_arbitration_removeIt = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      decode_arbitration_removeIt = 1'b1;
    end
  end

  assign decode_arbitration_flushIt = 1'b0;
  always @(*) begin
    decode_arbitration_flushNext = 1'b0;
    if(_zz_when) begin
      decode_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_haltItself = 1'b0;
    if(when_DBusSimplePlugin_l426) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_ShiftPlugins_l169) begin
      if(when_ShiftPlugins_l184) begin
        execute_arbitration_haltItself = 1'b1;
      end
    end
    if(when_CsrPlugin_l1180) begin
      if(execute_CsrPlugin_blockedBySideEffects) begin
        execute_arbitration_haltItself = 1'b1;
      end
    end
  end

  always @(*) begin
    execute_arbitration_haltByOther = 1'b0;
    if(when_DebugPlugin_l284) begin
      execute_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_removeIt = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_removeIt = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      execute_arbitration_removeIt = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_flushIt = 1'b0;
    if(when_DebugPlugin_l284) begin
      if(when_DebugPlugin_l287) begin
        execute_arbitration_flushIt = 1'b1;
      end
    end
  end

  always @(*) begin
    execute_arbitration_flushNext = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_flushNext = 1'b1;
    end
    if(when_DebugPlugin_l284) begin
      if(when_DebugPlugin_l287) begin
        execute_arbitration_flushNext = 1'b1;
      end
    end
  end

  always @(*) begin
    memory_arbitration_haltItself = 1'b0;
    if(when_DBusSimplePlugin_l479) begin
      memory_arbitration_haltItself = 1'b1;
    end
  end

  assign memory_arbitration_haltByOther = 1'b0;
  always @(*) begin
    memory_arbitration_removeIt = 1'b0;
    if(_zz_when_1) begin
      memory_arbitration_removeIt = 1'b1;
    end
    if(memory_arbitration_isFlushed) begin
      memory_arbitration_removeIt = 1'b1;
    end
  end

  assign memory_arbitration_flushIt = 1'b0;
  always @(*) begin
    memory_arbitration_flushNext = 1'b0;
    if(BranchPlugin_jumpInterface_valid) begin
      memory_arbitration_flushNext = 1'b1;
    end
    if(_zz_when_1) begin
      memory_arbitration_flushNext = 1'b1;
    end
  end

  assign writeBack_arbitration_haltItself = 1'b0;
  assign writeBack_arbitration_haltByOther = 1'b0;
  always @(*) begin
    writeBack_arbitration_removeIt = 1'b0;
    if(writeBack_arbitration_isFlushed) begin
      writeBack_arbitration_removeIt = 1'b1;
    end
  end

  assign writeBack_arbitration_flushIt = 1'b0;
  always @(*) begin
    writeBack_arbitration_flushNext = 1'b0;
    if(when_CsrPlugin_l1019) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(when_CsrPlugin_l1064) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
  end

  assign lastStageInstruction = writeBack_INSTRUCTION;
  assign lastStagePc = writeBack_PC;
  assign lastStageIsValid = writeBack_arbitration_isValid;
  assign lastStageIsFiring = writeBack_arbitration_isFiring;
  always @(*) begin
    IBusCachedPlugin_fetcherHalt = 1'b0;
    if(when_CsrPlugin_l922) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1019) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1064) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_DebugPlugin_l284) begin
      if(when_DebugPlugin_l287) begin
        IBusCachedPlugin_fetcherHalt = 1'b1;
      end
    end
    if(DebugPlugin_haltIt) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_DebugPlugin_l300) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_incomingInstruction = 1'b0;
    if(when_Fetcher_l240) begin
      IBusCachedPlugin_incomingInstruction = 1'b1;
    end
  end

  assign CsrPlugin_csrMapping_allowCsrSignal = 1'b0;
  assign CsrPlugin_csrMapping_readDataSignal = CsrPlugin_csrMapping_readDataInit;
  assign CsrPlugin_inWfi = 1'b0;
  always @(*) begin
    CsrPlugin_thirdPartyWake = 1'b0;
    if(DebugPlugin_haltIt) begin
      CsrPlugin_thirdPartyWake = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_valid = 1'b0;
    if(when_CsrPlugin_l1019) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
    if(when_CsrPlugin_l1064) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_CsrPlugin_l1019) begin
      CsrPlugin_jumpInterface_payload = {CsrPlugin_xtvec_base,2'b00};
    end
    if(when_CsrPlugin_l1064) begin
      case(switch_CsrPlugin_l1068)
        2'b11 : begin
          CsrPlugin_jumpInterface_payload = CsrPlugin_mepc;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CsrPlugin_forceMachineWire = 1'b0;
    if(DebugPlugin_godmode) begin
      CsrPlugin_forceMachineWire = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_allowInterrupts = 1'b1;
    if(when_DebugPlugin_l316) begin
      CsrPlugin_allowInterrupts = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_allowException = 1'b1;
    if(DebugPlugin_godmode) begin
      CsrPlugin_allowException = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_allowEbreakException = 1'b1;
    if(DebugPlugin_allowEBreak) begin
      CsrPlugin_allowEbreakException = 1'b0;
    end
  end

  assign IBusCachedPlugin_externalFlush = ({writeBack_arbitration_flushNext,{memory_arbitration_flushNext,{execute_arbitration_flushNext,decode_arbitration_flushNext}}} != 4'b0000);
  assign IBusCachedPlugin_jump_pcLoad_valid = ({CsrPlugin_jumpInterface_valid,BranchPlugin_jumpInterface_valid} != 2'b00);
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload = {BranchPlugin_jumpInterface_valid,CsrPlugin_jumpInterface_valid};
  assign IBusCachedPlugin_jump_pcLoad_payload = (_zz_IBusCachedPlugin_jump_pcLoad_payload_1[0] ? CsrPlugin_jumpInterface_payload : BranchPlugin_jumpInterface_payload);
  always @(*) begin
    IBusCachedPlugin_fetchPc_correction = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
  end

  assign IBusCachedPlugin_fetchPc_output_fire = (IBusCachedPlugin_fetchPc_output_valid && IBusCachedPlugin_fetchPc_output_ready);
  assign IBusCachedPlugin_fetchPc_corrected = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_correctionReg);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b0;
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b1;
    end
  end

  assign when_Fetcher_l131 = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_pcRegPropagate);
  assign IBusCachedPlugin_fetchPc_output_fire_1 = (IBusCachedPlugin_fetchPc_output_valid && IBusCachedPlugin_fetchPc_output_ready);
  assign when_Fetcher_l131_1 = ((! IBusCachedPlugin_fetchPc_output_valid) && IBusCachedPlugin_fetchPc_output_ready);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pc = (IBusCachedPlugin_fetchPc_pcReg + _zz_IBusCachedPlugin_fetchPc_pc);
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_fetchPc_redo_payload;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_jump_pcLoad_payload;
    end
    IBusCachedPlugin_fetchPc_pc[0] = 1'b0;
    IBusCachedPlugin_fetchPc_pc[1] = 1'b0;
  end

  always @(*) begin
    IBusCachedPlugin_fetchPc_flushed = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
  end

  assign when_Fetcher_l158 = (IBusCachedPlugin_fetchPc_booted && ((IBusCachedPlugin_fetchPc_output_ready || IBusCachedPlugin_fetchPc_correction) || IBusCachedPlugin_fetchPc_pcRegPropagate));
  assign IBusCachedPlugin_fetchPc_output_valid = ((! IBusCachedPlugin_fetcherHalt) && IBusCachedPlugin_fetchPc_booted);
  assign IBusCachedPlugin_fetchPc_output_payload = IBusCachedPlugin_fetchPc_pc;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_redoFetch = 1'b0;
    if(IBusCachedPlugin_rsp_redoFetch) begin
      IBusCachedPlugin_iBusRsp_redoFetch = 1'b1;
    end
  end

  assign IBusCachedPlugin_iBusRsp_stages_0_input_valid = IBusCachedPlugin_fetchPc_output_valid;
  assign IBusCachedPlugin_fetchPc_output_ready = IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_0_input_payload = IBusCachedPlugin_fetchPc_output_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b0;
    if(IBusCachedPlugin_cache_io_cpu_prefetch_haltIt) begin
      IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready = (! IBusCachedPlugin_iBusRsp_stages_0_halt);
  assign IBusCachedPlugin_iBusRsp_stages_0_input_ready = (IBusCachedPlugin_iBusRsp_stages_0_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_valid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_payload = IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b0;
    if(IBusCachedPlugin_mmuBus_busy) begin
      IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready = (! IBusCachedPlugin_iBusRsp_stages_1_halt);
  assign IBusCachedPlugin_iBusRsp_stages_1_input_ready = (IBusCachedPlugin_iBusRsp_stages_1_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_valid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_payload = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b0;
    if(when_IBusCachedPlugin_l267) begin
      IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready = (! IBusCachedPlugin_iBusRsp_stages_2_halt);
  assign IBusCachedPlugin_iBusRsp_stages_2_input_ready = (IBusCachedPlugin_iBusRsp_stages_2_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_valid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  assign IBusCachedPlugin_fetchPc_redo_valid = IBusCachedPlugin_iBusRsp_redoFetch;
  assign IBusCachedPlugin_fetchPc_redo_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  assign IBusCachedPlugin_iBusRsp_flush = ((decode_arbitration_removeIt || (decode_arbitration_flushNext && (! decode_arbitration_isStuck))) || IBusCachedPlugin_iBusRsp_redoFetch);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_ready = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready = ((1'b0 && (! _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1)) || IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1 = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_valid = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_payload = IBusCachedPlugin_fetchPc_pcReg;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_ready = ((1'b0 && (! IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid)) || IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_valid = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready = IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_payload = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_readyForError = 1'b1;
    if(when_Fetcher_l320) begin
      IBusCachedPlugin_iBusRsp_readyForError = 1'b0;
    end
  end

  assign when_Fetcher_l240 = (IBusCachedPlugin_iBusRsp_stages_1_input_valid || IBusCachedPlugin_iBusRsp_stages_2_input_valid);
  assign when_Fetcher_l320 = (! IBusCachedPlugin_pcValids_0);
  assign when_Fetcher_l329 = (! (! IBusCachedPlugin_iBusRsp_stages_1_input_ready));
  assign when_Fetcher_l329_1 = (! (! IBusCachedPlugin_iBusRsp_stages_2_input_ready));
  assign when_Fetcher_l329_2 = (! execute_arbitration_isStuck);
  assign when_Fetcher_l329_3 = (! memory_arbitration_isStuck);
  assign when_Fetcher_l329_4 = (! writeBack_arbitration_isStuck);
  assign IBusCachedPlugin_pcValids_0 = IBusCachedPlugin_injector_nextPcCalc_valids_1;
  assign IBusCachedPlugin_pcValids_1 = IBusCachedPlugin_injector_nextPcCalc_valids_2;
  assign IBusCachedPlugin_pcValids_2 = IBusCachedPlugin_injector_nextPcCalc_valids_3;
  assign IBusCachedPlugin_pcValids_3 = IBusCachedPlugin_injector_nextPcCalc_valids_4;
  assign IBusCachedPlugin_iBusRsp_output_ready = (! decode_arbitration_isStuck);
  always @(*) begin
    decode_arbitration_isValid = IBusCachedPlugin_iBusRsp_output_valid;
    case(switch_Fetcher_l362)
      3'b010 : begin
        decode_arbitration_isValid = 1'b1;
      end
      3'b011 : begin
        decode_arbitration_isValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign iBus_cmd_valid = IBusCachedPlugin_cache_io_mem_cmd_valid;
  always @(*) begin
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  end

  assign iBus_cmd_payload_size = IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  assign IBusCachedPlugin_s0_tightlyCoupledHit = 1'b0;
  assign IBusCachedPlugin_cache_io_cpu_prefetch_isValid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && (! IBusCachedPlugin_s0_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isValid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && (! IBusCachedPlugin_s1_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_isValid = IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  assign IBusCachedPlugin_mmuBus_cmd_0_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_virtualAddress = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  assign IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation = 1'b0;
  assign IBusCachedPlugin_mmuBus_end = (IBusCachedPlugin_iBusRsp_stages_1_input_ready || IBusCachedPlugin_externalFlush);
  assign IBusCachedPlugin_cache_io_cpu_decode_isValid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && (! IBusCachedPlugin_s2_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_decode_isStuck = (! IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_cache_io_cpu_decode_isUser = (CsrPlugin_privilege == 2'b00);
  assign IBusCachedPlugin_rsp_iBusRspOutputHalt = 1'b0;
  assign IBusCachedPlugin_rsp_issueDetected = 1'b0;
  always @(*) begin
    IBusCachedPlugin_rsp_redoFetch = 1'b0;
    if(when_IBusCachedPlugin_l239) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_cache_io_cpu_fill_valid = (IBusCachedPlugin_rsp_redoFetch && (! IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling));
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_cache_io_cpu_fill_valid = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_valid = 1'b0;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_payload_code = 4'bxxxx;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b1100;
    end
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b0001;
    end
  end

  assign IBusCachedPlugin_decodeExceptionPort_payload_badAddr = {IBusCachedPlugin_iBusRsp_stages_2_input_payload[31 : 2],2'b00};
  assign when_IBusCachedPlugin_l239 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling) && (! IBusCachedPlugin_rsp_issueDetected));
  assign when_IBusCachedPlugin_l244 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuException) && (! IBusCachedPlugin_rsp_issueDetected_1));
  assign when_IBusCachedPlugin_l250 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_cacheMiss) && (! IBusCachedPlugin_rsp_issueDetected_2));
  assign when_IBusCachedPlugin_l256 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_error) && (! IBusCachedPlugin_rsp_issueDetected_3));
  assign when_IBusCachedPlugin_l267 = (IBusCachedPlugin_rsp_issueDetected_4 || IBusCachedPlugin_rsp_iBusRspOutputHalt);
  assign IBusCachedPlugin_iBusRsp_output_valid = IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  assign IBusCachedPlugin_iBusRsp_stages_2_output_ready = IBusCachedPlugin_iBusRsp_output_ready;
  assign IBusCachedPlugin_iBusRsp_output_payload_rsp_inst = IBusCachedPlugin_cache_io_cpu_decode_data;
  assign IBusCachedPlugin_iBusRsp_output_payload_pc = IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  assign IBusCachedPlugin_cache_io_flush = (decode_arbitration_isValid && decode_FLUSH_ALL);
  assign _zz_dBus_cmd_valid = 1'b0;
  always @(*) begin
    execute_DBusSimplePlugin_skipCmd = 1'b0;
    if(execute_ALIGNEMENT_FAULT) begin
      execute_DBusSimplePlugin_skipCmd = 1'b1;
    end
  end

  assign dBus_cmd_valid = (((((execute_arbitration_isValid && execute_MEMORY_ENABLE) && (! execute_arbitration_isStuckByOthers)) && (! execute_arbitration_isFlushed)) && (! execute_DBusSimplePlugin_skipCmd)) && (! _zz_dBus_cmd_valid));
  assign dBus_cmd_payload_wr = execute_MEMORY_STORE;
  assign dBus_cmd_payload_size = execute_INSTRUCTION[13 : 12];
  always @(*) begin
    case(dBus_cmd_payload_size)
      2'b00 : begin
        _zz_dBus_cmd_payload_data = {{{execute_RS2[7 : 0],execute_RS2[7 : 0]},execute_RS2[7 : 0]},execute_RS2[7 : 0]};
      end
      2'b01 : begin
        _zz_dBus_cmd_payload_data = {execute_RS2[15 : 0],execute_RS2[15 : 0]};
      end
      default : begin
        _zz_dBus_cmd_payload_data = execute_RS2[31 : 0];
      end
    endcase
  end

  assign dBus_cmd_payload_data = _zz_dBus_cmd_payload_data;
  assign when_DBusSimplePlugin_l426 = ((((execute_arbitration_isValid && execute_MEMORY_ENABLE) && (! dBus_cmd_ready)) && (! execute_DBusSimplePlugin_skipCmd)) && (! _zz_dBus_cmd_valid));
  always @(*) begin
    case(dBus_cmd_payload_size)
      2'b00 : begin
        _zz_execute_DBusSimplePlugin_formalMask = 4'b0001;
      end
      2'b01 : begin
        _zz_execute_DBusSimplePlugin_formalMask = 4'b0011;
      end
      default : begin
        _zz_execute_DBusSimplePlugin_formalMask = 4'b1111;
      end
    endcase
  end

  assign execute_DBusSimplePlugin_formalMask = (_zz_execute_DBusSimplePlugin_formalMask <<< dBus_cmd_payload_address[1 : 0]);
  assign dBus_cmd_payload_address = execute_SRC_ADD;
  assign when_DBusSimplePlugin_l479 = (((memory_arbitration_isValid && memory_MEMORY_ENABLE) && (! memory_MEMORY_STORE)) && ((! dBus_rsp_ready) || 1'b0));
  always @(*) begin
    DBusSimplePlugin_memoryExceptionPort_valid = 1'b0;
    if(when_DBusSimplePlugin_l486) begin
      DBusSimplePlugin_memoryExceptionPort_valid = 1'b1;
    end
    if(memory_ALIGNEMENT_FAULT) begin
      DBusSimplePlugin_memoryExceptionPort_valid = 1'b1;
    end
    if(when_DBusSimplePlugin_l512) begin
      DBusSimplePlugin_memoryExceptionPort_valid = 1'b0;
    end
  end

  always @(*) begin
    DBusSimplePlugin_memoryExceptionPort_payload_code = 4'bxxxx;
    if(when_DBusSimplePlugin_l486) begin
      DBusSimplePlugin_memoryExceptionPort_payload_code = 4'b0101;
    end
    if(memory_ALIGNEMENT_FAULT) begin
      DBusSimplePlugin_memoryExceptionPort_payload_code = {1'd0, _zz_DBusSimplePlugin_memoryExceptionPort_payload_code};
    end
  end

  assign DBusSimplePlugin_memoryExceptionPort_payload_badAddr = memory_REGFILE_WRITE_DATA;
  assign when_DBusSimplePlugin_l486 = ((dBus_rsp_ready && dBus_rsp_error) && (! memory_MEMORY_STORE));
  assign when_DBusSimplePlugin_l512 = (! ((memory_arbitration_isValid && memory_MEMORY_ENABLE) && (1'b1 || (! memory_arbitration_isStuckByOthers))));
  always @(*) begin
    writeBack_DBusSimplePlugin_rspShifted = writeBack_MEMORY_READ_DATA;
    case(writeBack_MEMORY_ADDRESS_LOW)
      2'b01 : begin
        writeBack_DBusSimplePlugin_rspShifted[7 : 0] = writeBack_MEMORY_READ_DATA[15 : 8];
      end
      2'b10 : begin
        writeBack_DBusSimplePlugin_rspShifted[15 : 0] = writeBack_MEMORY_READ_DATA[31 : 16];
      end
      2'b11 : begin
        writeBack_DBusSimplePlugin_rspShifted[7 : 0] = writeBack_MEMORY_READ_DATA[31 : 24];
      end
      default : begin
      end
    endcase
  end

  assign switch_Misc_l200 = writeBack_INSTRUCTION[13 : 12];
  assign _zz_writeBack_DBusSimplePlugin_rspFormated = (writeBack_DBusSimplePlugin_rspShifted[7] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[31] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[30] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[29] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[28] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[27] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[26] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[25] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[24] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[23] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[22] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[21] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[20] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[19] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[18] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[17] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[16] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[15] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[14] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[13] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[12] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[11] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[10] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[9] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[8] = _zz_writeBack_DBusSimplePlugin_rspFormated;
    _zz_writeBack_DBusSimplePlugin_rspFormated_1[7 : 0] = writeBack_DBusSimplePlugin_rspShifted[7 : 0];
  end

  assign _zz_writeBack_DBusSimplePlugin_rspFormated_2 = (writeBack_DBusSimplePlugin_rspShifted[15] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[31] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[30] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[29] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[28] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[27] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[26] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[25] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[24] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[23] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[22] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[21] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[20] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[19] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[18] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[17] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[16] = _zz_writeBack_DBusSimplePlugin_rspFormated_2;
    _zz_writeBack_DBusSimplePlugin_rspFormated_3[15 : 0] = writeBack_DBusSimplePlugin_rspShifted[15 : 0];
  end

  always @(*) begin
    case(switch_Misc_l200)
      2'b00 : begin
        writeBack_DBusSimplePlugin_rspFormated = _zz_writeBack_DBusSimplePlugin_rspFormated_1;
      end
      2'b01 : begin
        writeBack_DBusSimplePlugin_rspFormated = _zz_writeBack_DBusSimplePlugin_rspFormated_3;
      end
      default : begin
        writeBack_DBusSimplePlugin_rspFormated = writeBack_DBusSimplePlugin_rspShifted;
      end
    endcase
  end

  assign when_DBusSimplePlugin_l558 = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
  assign IBusCachedPlugin_mmuBus_rsp_physicalAddress = IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  assign IBusCachedPlugin_mmuBus_rsp_allowRead = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_allowWrite = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_allowExecute = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_isIoAccess = IBusCachedPlugin_mmuBus_rsp_physicalAddress[31];
  assign IBusCachedPlugin_mmuBus_rsp_isPaging = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_exception = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_refilling = 1'b0;
  assign IBusCachedPlugin_mmuBus_busy = 1'b0;
  assign _zz_decode_ENV_CTRL_3 = ((decode_INSTRUCTION & 32'h00004050) == 32'h00004050);
  assign _zz_decode_ENV_CTRL_4 = ((decode_INSTRUCTION & 32'h00000004) == 32'h00000004);
  assign _zz_decode_ENV_CTRL_5 = ((decode_INSTRUCTION & 32'h00000050) == 32'h00000010);
  assign _zz_decode_ENV_CTRL_6 = ((decode_INSTRUCTION & 32'h00000048) == 32'h00000048);
  assign _zz_decode_ENV_CTRL_2 = {(((decode_INSTRUCTION & _zz__zz_decode_ENV_CTRL_2) == 32'h00100050) != 1'b0),{((_zz__zz_decode_ENV_CTRL_2_1 == _zz__zz_decode_ENV_CTRL_2_2) != 1'b0),{(_zz__zz_decode_ENV_CTRL_2_3 != 1'b0),{(_zz__zz_decode_ENV_CTRL_2_4 != _zz__zz_decode_ENV_CTRL_2_9),{_zz__zz_decode_ENV_CTRL_2_10,{_zz__zz_decode_ENV_CTRL_2_12,_zz__zz_decode_ENV_CTRL_2_14}}}}}};
  assign _zz_decode_SRC1_CTRL_2 = _zz_decode_ENV_CTRL_2[2 : 1];
  assign _zz_decode_SRC1_CTRL_1 = _zz_decode_SRC1_CTRL_2;
  assign _zz_decode_ALU_CTRL_2 = _zz_decode_ENV_CTRL_2[7 : 6];
  assign _zz_decode_ALU_CTRL_1 = _zz_decode_ALU_CTRL_2;
  assign _zz_decode_SRC2_CTRL_2 = _zz_decode_ENV_CTRL_2[9 : 8];
  assign _zz_decode_SRC2_CTRL_1 = _zz_decode_SRC2_CTRL_2;
  assign _zz_decode_ALU_BITWISE_CTRL_2 = _zz_decode_ENV_CTRL_2[18 : 17];
  assign _zz_decode_ALU_BITWISE_CTRL_1 = _zz_decode_ALU_BITWISE_CTRL_2;
  assign _zz_decode_SHIFT_CTRL_2 = _zz_decode_ENV_CTRL_2[21 : 20];
  assign _zz_decode_SHIFT_CTRL_1 = _zz_decode_SHIFT_CTRL_2;
  assign _zz_decode_BRANCH_CTRL_2 = _zz_decode_ENV_CTRL_2[23 : 22];
  assign _zz_decode_BRANCH_CTRL_1 = _zz_decode_BRANCH_CTRL_2;
  assign _zz_decode_ENV_CTRL_7 = _zz_decode_ENV_CTRL_2[26 : 25];
  assign _zz_decode_ENV_CTRL_1 = _zz_decode_ENV_CTRL_7;
  assign decodeExceptionPort_valid = (decode_arbitration_isValid && (! decode_LEGAL_INSTRUCTION));
  assign decodeExceptionPort_payload_code = 4'b0010;
  assign decodeExceptionPort_payload_badAddr = decode_INSTRUCTION;
  assign when_RegFilePlugin_l63 = (decode_INSTRUCTION[11 : 7] == 5'h0);
  assign decode_RegFilePlugin_regFileReadAddress1 = decode_INSTRUCTION_ANTICIPATED[19 : 15];
  assign decode_RegFilePlugin_regFileReadAddress2 = decode_INSTRUCTION_ANTICIPATED[24 : 20];
  assign decode_RegFilePlugin_rs1Data = _zz_RegFilePlugin_regFile_port0;
  assign decode_RegFilePlugin_rs2Data = _zz_RegFilePlugin_regFile_port1;
  always @(*) begin
    lastStageRegFileWrite_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
    if(_zz_2) begin
      lastStageRegFileWrite_valid = 1'b1;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
    if(_zz_2) begin
      lastStageRegFileWrite_payload_address = 5'h0;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_data = _zz_lastStageRegFileWrite_payload_data;
    if(_zz_2) begin
      lastStageRegFileWrite_payload_data = 32'h0;
    end
  end

  always @(*) begin
    case(execute_ALU_BITWISE_CTRL)
      2'b10 : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 & execute_SRC2);
      end
      2'b01 : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 | execute_SRC2);
      end
      default : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 ^ execute_SRC2);
      end
    endcase
  end

  always @(*) begin
    case(execute_ALU_CTRL)
      2'b10 : begin
        _zz_execute_REGFILE_WRITE_DATA = execute_IntAluPlugin_bitwise;
      end
      2'b01 : begin
        _zz_execute_REGFILE_WRITE_DATA = {31'd0, _zz__zz_execute_REGFILE_WRITE_DATA};
      end
      default : begin
        _zz_execute_REGFILE_WRITE_DATA = execute_SRC_ADD_SUB;
      end
    endcase
  end

  always @(*) begin
    case(execute_SRC1_CTRL)
      2'b00 : begin
        _zz_execute_SRC1 = execute_RS1;
      end
      2'b10 : begin
        _zz_execute_SRC1 = {29'd0, _zz__zz_execute_SRC1};
      end
      2'b01 : begin
        _zz_execute_SRC1 = {execute_INSTRUCTION[31 : 12],12'h0};
      end
      default : begin
        _zz_execute_SRC1 = {27'd0, _zz__zz_execute_SRC1_1};
      end
    endcase
  end

  assign _zz_execute_SRC2_1 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_SRC2_2[19] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[18] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[17] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[16] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[15] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[14] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[13] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[12] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[11] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[10] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[9] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[8] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[7] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[6] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[5] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[4] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[3] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[2] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[1] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[0] = _zz_execute_SRC2_1;
  end

  assign _zz_execute_SRC2_3 = _zz__zz_execute_SRC2_3[11];
  always @(*) begin
    _zz_execute_SRC2_4[19] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[18] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[17] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[16] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[15] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[14] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[13] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[12] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[11] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[10] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[9] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[8] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[7] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[6] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[5] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[4] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[3] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[2] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[1] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[0] = _zz_execute_SRC2_3;
  end

  always @(*) begin
    case(execute_SRC2_CTRL)
      2'b00 : begin
        _zz_execute_SRC2_5 = execute_RS2;
      end
      2'b01 : begin
        _zz_execute_SRC2_5 = {_zz_execute_SRC2_2,execute_INSTRUCTION[31 : 20]};
      end
      2'b10 : begin
        _zz_execute_SRC2_5 = {_zz_execute_SRC2_4,{execute_INSTRUCTION[31 : 25],execute_INSTRUCTION[11 : 7]}};
      end
      default : begin
        _zz_execute_SRC2_5 = _zz_execute_SRC2;
      end
    endcase
  end

  always @(*) begin
    execute_SrcPlugin_addSub = _zz_execute_SrcPlugin_addSub;
    if(execute_SRC2_FORCE_ZERO) begin
      execute_SrcPlugin_addSub = execute_SRC1;
    end
  end

  assign execute_SrcPlugin_less = ((execute_SRC1[31] == execute_SRC2[31]) ? execute_SrcPlugin_addSub[31] : (execute_SRC_LESS_UNSIGNED ? execute_SRC2[31] : execute_SRC1[31]));
  assign execute_LightShifterPlugin_isShift = (execute_SHIFT_CTRL != 2'b00);
  assign execute_LightShifterPlugin_amplitude = (execute_LightShifterPlugin_isActive ? execute_LightShifterPlugin_amplitudeReg : execute_SRC2[4 : 0]);
  assign execute_LightShifterPlugin_shiftInput = (execute_LightShifterPlugin_isActive ? memory_REGFILE_WRITE_DATA : execute_SRC1);
  assign execute_LightShifterPlugin_done = (execute_LightShifterPlugin_amplitude[4 : 1] == 4'b0000);
  assign when_ShiftPlugins_l169 = ((execute_arbitration_isValid && execute_LightShifterPlugin_isShift) && (execute_SRC2[4 : 0] != 5'h0));
  always @(*) begin
    case(execute_SHIFT_CTRL)
      2'b01 : begin
        _zz_execute_to_memory_REGFILE_WRITE_DATA_1 = (execute_LightShifterPlugin_shiftInput <<< 1);
      end
      default : begin
        _zz_execute_to_memory_REGFILE_WRITE_DATA_1 = _zz__zz_execute_to_memory_REGFILE_WRITE_DATA_1;
      end
    endcase
  end

  assign when_ShiftPlugins_l175 = (! execute_arbitration_isStuckByOthers);
  assign when_ShiftPlugins_l184 = (! execute_LightShifterPlugin_done);
  always @(*) begin
    HazardSimplePlugin_src0Hazard = 1'b0;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr0Match) begin
        HazardSimplePlugin_src0Hazard = 1'b1;
      end
    end
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l59) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l59_1) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l59_2) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l105) begin
      HazardSimplePlugin_src0Hazard = 1'b0;
    end
  end

  always @(*) begin
    HazardSimplePlugin_src1Hazard = 1'b0;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr1Match) begin
        HazardSimplePlugin_src1Hazard = 1'b1;
      end
    end
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l62) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l62_1) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l62_2) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l108) begin
      HazardSimplePlugin_src1Hazard = 1'b0;
    end
  end

  assign HazardSimplePlugin_writeBackWrites_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
  assign HazardSimplePlugin_writeBackWrites_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
  assign HazardSimplePlugin_writeBackWrites_payload_data = _zz_lastStageRegFileWrite_payload_data;
  assign HazardSimplePlugin_addr0Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[19 : 15]);
  assign HazardSimplePlugin_addr1Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l59 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l62 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l57 = (writeBack_arbitration_isValid && writeBack_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58 = (1'b1 || (! 1'b1));
  assign when_HazardSimplePlugin_l59_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l62_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l57_1 = (memory_arbitration_isValid && memory_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_1 = (1'b1 || (! memory_BYPASSABLE_MEMORY_STAGE));
  assign when_HazardSimplePlugin_l59_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l62_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l57_2 = (execute_arbitration_isValid && execute_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_2 = (1'b1 || (! execute_BYPASSABLE_EXECUTE_STAGE));
  assign when_HazardSimplePlugin_l105 = (! decode_RS1_USE);
  assign when_HazardSimplePlugin_l108 = (! decode_RS2_USE);
  assign when_HazardSimplePlugin_l113 = (decode_arbitration_isValid && (HazardSimplePlugin_src0Hazard || HazardSimplePlugin_src1Hazard));
  assign execute_BranchPlugin_eq = (execute_SRC1 == execute_SRC2);
  assign switch_Misc_l200_1 = execute_INSTRUCTION[14 : 12];
  always @(*) begin
    casez(switch_Misc_l200_1)
      3'b000 : begin
        _zz_execute_BRANCH_DO = execute_BranchPlugin_eq;
      end
      3'b001 : begin
        _zz_execute_BRANCH_DO = (! execute_BranchPlugin_eq);
      end
      3'b1?1 : begin
        _zz_execute_BRANCH_DO = (! execute_SRC_LESS);
      end
      default : begin
        _zz_execute_BRANCH_DO = execute_SRC_LESS;
      end
    endcase
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      2'b00 : begin
        _zz_execute_BRANCH_DO_1 = 1'b0;
      end
      2'b10 : begin
        _zz_execute_BRANCH_DO_1 = 1'b1;
      end
      2'b11 : begin
        _zz_execute_BRANCH_DO_1 = 1'b1;
      end
      default : begin
        _zz_execute_BRANCH_DO_1 = _zz_execute_BRANCH_DO;
      end
    endcase
  end

  assign execute_BranchPlugin_branch_src1 = ((execute_BRANCH_CTRL == 2'b11) ? execute_RS1 : execute_PC);
  assign _zz_execute_BranchPlugin_branch_src2 = _zz__zz_execute_BranchPlugin_branch_src2[19];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_1[10] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[9] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[8] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[7] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[6] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[5] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[4] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[3] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[2] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[1] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[0] = _zz_execute_BranchPlugin_branch_src2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_2 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_3[19] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[18] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[17] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[16] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[15] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[14] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[13] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[12] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[11] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[10] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[9] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[8] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[7] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[6] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[5] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[4] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[3] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[2] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[1] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[0] = _zz_execute_BranchPlugin_branch_src2_2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_4 = _zz__zz_execute_BranchPlugin_branch_src2_4[11];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_5[18] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[17] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[16] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[15] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[14] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[13] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[12] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[11] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[10] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[9] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[8] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[7] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[6] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[5] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[4] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[3] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[2] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[1] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[0] = _zz_execute_BranchPlugin_branch_src2_4;
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      2'b10 : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {{_zz_execute_BranchPlugin_branch_src2_1,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]}},1'b0};
      end
      2'b11 : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {_zz_execute_BranchPlugin_branch_src2_3,execute_INSTRUCTION[31 : 20]};
      end
      default : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {{_zz_execute_BranchPlugin_branch_src2_5,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]}},1'b0};
      end
    endcase
  end

  assign execute_BranchPlugin_branch_src2 = _zz_execute_BranchPlugin_branch_src2_6;
  assign execute_BranchPlugin_branchAdder = (execute_BranchPlugin_branch_src1 + execute_BranchPlugin_branch_src2);
  assign BranchPlugin_jumpInterface_valid = ((memory_arbitration_isValid && memory_BRANCH_DO) && (! 1'b0));
  assign BranchPlugin_jumpInterface_payload = memory_BRANCH_CALC;
  assign BranchPlugin_branchExceptionPort_valid = ((memory_arbitration_isValid && memory_BRANCH_DO) && BranchPlugin_jumpInterface_payload[1]);
  assign BranchPlugin_branchExceptionPort_payload_code = 4'b0000;
  assign BranchPlugin_branchExceptionPort_payload_badAddr = BranchPlugin_jumpInterface_payload;
  always @(*) begin
    CsrPlugin_privilege = 2'b11;
    if(CsrPlugin_forceMachineWire) begin
      CsrPlugin_privilege = 2'b11;
    end
  end

  assign CsrPlugin_misa_base = 2'b01;
  assign CsrPlugin_misa_extensions = 26'h0000042;
  assign _zz_when_CsrPlugin_l952 = (CsrPlugin_mip_MTIP && CsrPlugin_mie_MTIE);
  assign _zz_when_CsrPlugin_l952_1 = (CsrPlugin_mip_MSIP && CsrPlugin_mie_MSIE);
  assign _zz_when_CsrPlugin_l952_2 = (CsrPlugin_mip_MEIP && CsrPlugin_mie_MEIE);
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped = 2'b11;
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege = ((CsrPlugin_privilege < CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped) ? CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped : CsrPlugin_privilege);
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code = {decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid};
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1[0];
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_2 = {BranchPlugin_branchExceptionPort_valid,DBusSimplePlugin_memoryExceptionPort_valid};
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3 = _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3[0];
  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_decode = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_execute = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_memory = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
    if(_zz_when_1) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory = 1'b1;
    end
    if(memory_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
    if(writeBack_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = 1'b0;
    end
  end

  assign when_CsrPlugin_l909 = (! decode_arbitration_isStuck);
  assign when_CsrPlugin_l909_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l909_2 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l909_3 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l922 = ({CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValids_memory,{CsrPlugin_exceptionPortCtrl_exceptionValids_execute,CsrPlugin_exceptionPortCtrl_exceptionValids_decode}}} != 4'b0000);
  assign CsrPlugin_exceptionPendings_0 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  assign CsrPlugin_exceptionPendings_1 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  assign CsrPlugin_exceptionPendings_2 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  assign CsrPlugin_exceptionPendings_3 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  assign when_CsrPlugin_l946 = (CsrPlugin_mstatus_MIE || (CsrPlugin_privilege < 2'b11));
  assign when_CsrPlugin_l952 = ((_zz_when_CsrPlugin_l952 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l952_1 = ((_zz_when_CsrPlugin_l952_1 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l952_2 = ((_zz_when_CsrPlugin_l952_2 && 1'b1) && (! 1'b0));
  assign CsrPlugin_exception = (CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack && CsrPlugin_allowException);
  assign CsrPlugin_lastStageWasWfi = 1'b0;
  assign CsrPlugin_pipelineLiberator_active = ((CsrPlugin_interrupt_valid && CsrPlugin_allowInterrupts) && decode_arbitration_isValid);
  assign when_CsrPlugin_l980 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l980_1 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l980_2 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l985 = ((! CsrPlugin_pipelineLiberator_active) || decode_arbitration_removeIt);
  always @(*) begin
    CsrPlugin_pipelineLiberator_done = CsrPlugin_pipelineLiberator_pcValids_2;
    if(when_CsrPlugin_l991) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
    if(CsrPlugin_hadException) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
  end

  assign when_CsrPlugin_l991 = ({CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory,CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute}} != 3'b000);
  assign CsrPlugin_interruptJump = ((CsrPlugin_interrupt_valid && CsrPlugin_pipelineLiberator_done) && CsrPlugin_allowInterrupts);
  always @(*) begin
    CsrPlugin_targetPrivilege = CsrPlugin_interrupt_targetPrivilege;
    if(CsrPlugin_hadException) begin
      CsrPlugin_targetPrivilege = CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
    end
  end

  always @(*) begin
    CsrPlugin_trapCause = CsrPlugin_interrupt_code;
    if(CsrPlugin_hadException) begin
      CsrPlugin_trapCause = CsrPlugin_exceptionPortCtrl_exceptionContext_code;
    end
  end

  always @(*) begin
    CsrPlugin_xtvec_mode = 2'bxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_mode = CsrPlugin_mtvec_mode;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_xtvec_base = 30'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_base = CsrPlugin_mtvec_base;
      end
      default : begin
      end
    endcase
  end

  assign when_CsrPlugin_l1019 = (CsrPlugin_hadException || CsrPlugin_interruptJump);
  assign when_CsrPlugin_l1064 = (writeBack_arbitration_isValid && (writeBack_ENV_CTRL == 2'b01));
  assign switch_CsrPlugin_l1068 = writeBack_INSTRUCTION[29 : 28];
  assign contextSwitching = CsrPlugin_jumpInterface_valid;
  assign when_CsrPlugin_l1116 = ({(writeBack_arbitration_isValid && (writeBack_ENV_CTRL == 2'b01)),{(memory_arbitration_isValid && (memory_ENV_CTRL == 2'b01)),(execute_arbitration_isValid && (execute_ENV_CTRL == 2'b01))}} != 3'b000);
  assign execute_CsrPlugin_blockedBySideEffects = (({writeBack_arbitration_isValid,memory_arbitration_isValid} != 2'b00) || 1'b0);
  always @(*) begin
    execute_CsrPlugin_illegalAccess = 1'b1;
    if(execute_CsrPlugin_csr_768) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_836) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_772) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_773) begin
      if(execute_CSR_WRITE_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_833) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_834) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_835) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3008) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_4032) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(CsrPlugin_csrMapping_allowCsrSignal) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(when_CsrPlugin_l1297) begin
      execute_CsrPlugin_illegalAccess = 1'b1;
    end
    if(when_CsrPlugin_l1302) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_illegalInstruction = 1'b0;
    if(when_CsrPlugin_l1136) begin
      if(when_CsrPlugin_l1137) begin
        execute_CsrPlugin_illegalInstruction = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrPlugin_selfException_valid = 1'b0;
    if(when_CsrPlugin_l1144) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_selfException_payload_code = 4'bxxxx;
    if(when_CsrPlugin_l1144) begin
      case(CsrPlugin_privilege)
        2'b00 : begin
          CsrPlugin_selfException_payload_code = 4'b1000;
        end
        default : begin
          CsrPlugin_selfException_payload_code = 4'b1011;
        end
      endcase
    end
  end

  assign CsrPlugin_selfException_payload_badAddr = execute_INSTRUCTION;
  assign when_CsrPlugin_l1136 = (execute_arbitration_isValid && (execute_ENV_CTRL == 2'b01));
  assign when_CsrPlugin_l1137 = (CsrPlugin_privilege < execute_INSTRUCTION[29 : 28]);
  assign when_CsrPlugin_l1144 = (execute_arbitration_isValid && (execute_ENV_CTRL == 2'b10));
  always @(*) begin
    execute_CsrPlugin_writeInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_WRITE_OPCODE);
    if(when_CsrPlugin_l1297) begin
      execute_CsrPlugin_writeInstruction = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_readInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_READ_OPCODE);
    if(when_CsrPlugin_l1297) begin
      execute_CsrPlugin_readInstruction = 1'b0;
    end
  end

  assign execute_CsrPlugin_writeEnable = (execute_CsrPlugin_writeInstruction && (! execute_arbitration_isStuck));
  assign execute_CsrPlugin_readEnable = (execute_CsrPlugin_readInstruction && (! execute_arbitration_isStuck));
  assign CsrPlugin_csrMapping_hazardFree = (! execute_CsrPlugin_blockedBySideEffects);
  assign execute_CsrPlugin_readToWriteData = CsrPlugin_csrMapping_readDataSignal;
  assign switch_Misc_l200_2 = execute_INSTRUCTION[13];
  always @(*) begin
    case(switch_Misc_l200_2)
      1'b0 : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = execute_SRC1;
      end
      default : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = (execute_INSTRUCTION[12] ? (execute_CsrPlugin_readToWriteData & (~ execute_SRC1)) : (execute_CsrPlugin_readToWriteData | execute_SRC1));
      end
    endcase
  end

  assign CsrPlugin_csrMapping_writeDataSignal = _zz_CsrPlugin_csrMapping_writeDataSignal;
  assign when_CsrPlugin_l1176 = (execute_arbitration_isValid && execute_IS_CSR);
  assign when_CsrPlugin_l1180 = (execute_arbitration_isValid && (execute_IS_CSR || 1'b0));
  assign execute_CsrPlugin_csrAddress = execute_INSTRUCTION[31 : 20];
  assign _zz_CsrPlugin_csrMapping_readDataInit_1 = (_zz_CsrPlugin_csrMapping_readDataInit & externalInterruptArray_regNext);
  assign externalInterrupt = (_zz_CsrPlugin_csrMapping_readDataInit_1 != 32'h0);
  assign when_DebugPlugin_l225 = (DebugPlugin_haltIt && (! DebugPlugin_isPipBusy));
  assign DebugPlugin_allowEBreak = (DebugPlugin_debugUsed && (! DebugPlugin_disableEbreak));
  always @(*) begin
    debug_bus_cmd_ready = 1'b1;
    if(debug_bus_cmd_valid) begin
      case(switch_DebugPlugin_l256)
        6'h01 : begin
          if(debug_bus_cmd_payload_wr) begin
            debug_bus_cmd_ready = IBusCachedPlugin_injectionPort_ready;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    debug_bus_rsp_data = DebugPlugin_busReadDataReg;
    if(when_DebugPlugin_l244) begin
      debug_bus_rsp_data[0] = DebugPlugin_resetIt;
      debug_bus_rsp_data[1] = DebugPlugin_haltIt;
      debug_bus_rsp_data[2] = DebugPlugin_isPipBusy;
      debug_bus_rsp_data[3] = DebugPlugin_haltedByBreak;
      debug_bus_rsp_data[4] = DebugPlugin_stepIt;
    end
  end

  assign when_DebugPlugin_l244 = (! _zz_when_DebugPlugin_l244);
  always @(*) begin
    IBusCachedPlugin_injectionPort_valid = 1'b0;
    if(debug_bus_cmd_valid) begin
      case(switch_DebugPlugin_l256)
        6'h01 : begin
          if(debug_bus_cmd_payload_wr) begin
            IBusCachedPlugin_injectionPort_valid = 1'b1;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign IBusCachedPlugin_injectionPort_payload = debug_bus_cmd_payload_data;
  assign switch_DebugPlugin_l256 = debug_bus_cmd_payload_address[7 : 2];
  assign when_DebugPlugin_l260 = debug_bus_cmd_payload_data[16];
  assign when_DebugPlugin_l260_1 = debug_bus_cmd_payload_data[24];
  assign when_DebugPlugin_l261 = debug_bus_cmd_payload_data[17];
  assign when_DebugPlugin_l261_1 = debug_bus_cmd_payload_data[25];
  assign when_DebugPlugin_l262 = debug_bus_cmd_payload_data[25];
  assign when_DebugPlugin_l263 = debug_bus_cmd_payload_data[25];
  assign when_DebugPlugin_l264 = debug_bus_cmd_payload_data[18];
  assign when_DebugPlugin_l264_1 = debug_bus_cmd_payload_data[26];
  assign when_DebugPlugin_l284 = (execute_arbitration_isValid && execute_DO_EBREAK);
  assign when_DebugPlugin_l287 = (({writeBack_arbitration_isValid,memory_arbitration_isValid} != 2'b00) == 1'b0);
  assign when_DebugPlugin_l300 = (DebugPlugin_stepIt && IBusCachedPlugin_incomingInstruction);
  assign debug_resetOut = DebugPlugin_resetIt_regNext;
  assign when_DebugPlugin_l316 = (DebugPlugin_haltIt || DebugPlugin_stepIt);
  assign when_Pipeline_l124 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_1 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_2 = ((! writeBack_arbitration_isStuck) && (! CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack));
  assign when_Pipeline_l124_3 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_4 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_5 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_6 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_7 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_8 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_SRC1_CTRL_1 = decode_SRC1_CTRL;
  assign _zz_decode_SRC1_CTRL = _zz_decode_SRC1_CTRL_1;
  assign when_Pipeline_l124_9 = (! execute_arbitration_isStuck);
  assign _zz_execute_SRC1_CTRL = decode_to_execute_SRC1_CTRL;
  assign when_Pipeline_l124_10 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_11 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_12 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_13 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_ALU_CTRL_1 = decode_ALU_CTRL;
  assign _zz_decode_ALU_CTRL = _zz_decode_ALU_CTRL_1;
  assign when_Pipeline_l124_14 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_CTRL = decode_to_execute_ALU_CTRL;
  assign _zz_decode_to_execute_SRC2_CTRL_1 = decode_SRC2_CTRL;
  assign _zz_decode_SRC2_CTRL = _zz_decode_SRC2_CTRL_1;
  assign when_Pipeline_l124_15 = (! execute_arbitration_isStuck);
  assign _zz_execute_SRC2_CTRL = decode_to_execute_SRC2_CTRL;
  assign when_Pipeline_l124_16 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_17 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_18 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_19 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_20 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_21 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_22 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_23 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_24 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_25 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL_1 = decode_ALU_BITWISE_CTRL;
  assign _zz_decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL_1;
  assign when_Pipeline_l124_26 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_BITWISE_CTRL = decode_to_execute_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL_1 = decode_SHIFT_CTRL;
  assign _zz_decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL_1;
  assign when_Pipeline_l124_27 = (! execute_arbitration_isStuck);
  assign _zz_execute_SHIFT_CTRL = decode_to_execute_SHIFT_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL_1 = decode_BRANCH_CTRL;
  assign _zz_decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL_1;
  assign when_Pipeline_l124_28 = (! execute_arbitration_isStuck);
  assign _zz_execute_BRANCH_CTRL = decode_to_execute_BRANCH_CTRL;
  assign when_Pipeline_l124_29 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_ENV_CTRL_1 = decode_ENV_CTRL;
  assign _zz_execute_to_memory_ENV_CTRL_1 = execute_ENV_CTRL;
  assign _zz_memory_to_writeBack_ENV_CTRL_1 = memory_ENV_CTRL;
  assign _zz_decode_ENV_CTRL = _zz_decode_ENV_CTRL_1;
  assign when_Pipeline_l124_30 = (! execute_arbitration_isStuck);
  assign _zz_execute_ENV_CTRL = decode_to_execute_ENV_CTRL;
  assign when_Pipeline_l124_31 = (! memory_arbitration_isStuck);
  assign _zz_memory_ENV_CTRL = execute_to_memory_ENV_CTRL;
  assign when_Pipeline_l124_32 = (! writeBack_arbitration_isStuck);
  assign _zz_writeBack_ENV_CTRL = memory_to_writeBack_ENV_CTRL;
  assign when_Pipeline_l124_33 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_34 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_35 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_36 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_37 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_38 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_39 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_40 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_41 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_42 = ((! memory_arbitration_isStuck) && (! execute_arbitration_isStuckByOthers));
  assign when_Pipeline_l124_43 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_44 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_45 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_46 = (! writeBack_arbitration_isStuck);
  assign decode_arbitration_isFlushed = (({writeBack_arbitration_flushNext,{memory_arbitration_flushNext,execute_arbitration_flushNext}} != 3'b000) || ({writeBack_arbitration_flushIt,{memory_arbitration_flushIt,{execute_arbitration_flushIt,decode_arbitration_flushIt}}} != 4'b0000));
  assign execute_arbitration_isFlushed = (({writeBack_arbitration_flushNext,memory_arbitration_flushNext} != 2'b00) || ({writeBack_arbitration_flushIt,{memory_arbitration_flushIt,execute_arbitration_flushIt}} != 3'b000));
  assign memory_arbitration_isFlushed = ((writeBack_arbitration_flushNext != 1'b0) || ({writeBack_arbitration_flushIt,memory_arbitration_flushIt} != 2'b00));
  assign writeBack_arbitration_isFlushed = (1'b0 || (writeBack_arbitration_flushIt != 1'b0));
  assign decode_arbitration_isStuckByOthers = (decode_arbitration_haltByOther || (((1'b0 || execute_arbitration_isStuck) || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign decode_arbitration_isStuck = (decode_arbitration_haltItself || decode_arbitration_isStuckByOthers);
  assign decode_arbitration_isMoving = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign decode_arbitration_isFiring = ((decode_arbitration_isValid && (! decode_arbitration_isStuck)) && (! decode_arbitration_removeIt));
  assign execute_arbitration_isStuckByOthers = (execute_arbitration_haltByOther || ((1'b0 || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign execute_arbitration_isStuck = (execute_arbitration_haltItself || execute_arbitration_isStuckByOthers);
  assign execute_arbitration_isMoving = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign execute_arbitration_isFiring = ((execute_arbitration_isValid && (! execute_arbitration_isStuck)) && (! execute_arbitration_removeIt));
  assign memory_arbitration_isStuckByOthers = (memory_arbitration_haltByOther || (1'b0 || writeBack_arbitration_isStuck));
  assign memory_arbitration_isStuck = (memory_arbitration_haltItself || memory_arbitration_isStuckByOthers);
  assign memory_arbitration_isMoving = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  assign memory_arbitration_isFiring = ((memory_arbitration_isValid && (! memory_arbitration_isStuck)) && (! memory_arbitration_removeIt));
  assign writeBack_arbitration_isStuckByOthers = (writeBack_arbitration_haltByOther || 1'b0);
  assign writeBack_arbitration_isStuck = (writeBack_arbitration_haltItself || writeBack_arbitration_isStuckByOthers);
  assign writeBack_arbitration_isMoving = ((! writeBack_arbitration_isStuck) && (! writeBack_arbitration_removeIt));
  assign writeBack_arbitration_isFiring = ((writeBack_arbitration_isValid && (! writeBack_arbitration_isStuck)) && (! writeBack_arbitration_removeIt));
  assign when_Pipeline_l151 = ((! execute_arbitration_isStuck) || execute_arbitration_removeIt);
  assign when_Pipeline_l154 = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign when_Pipeline_l151_1 = ((! memory_arbitration_isStuck) || memory_arbitration_removeIt);
  assign when_Pipeline_l154_1 = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign when_Pipeline_l151_2 = ((! writeBack_arbitration_isStuck) || writeBack_arbitration_removeIt);
  assign when_Pipeline_l154_2 = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  always @(*) begin
    IBusCachedPlugin_injectionPort_ready = 1'b0;
    case(switch_Fetcher_l362)
      3'b100 : begin
        IBusCachedPlugin_injectionPort_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign when_Fetcher_l378 = (! decode_arbitration_isStuck);
  assign when_CsrPlugin_l1264 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_2 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_3 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_4 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_5 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_6 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_7 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1264_8 = (! execute_arbitration_isStuck);
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_2 = 32'h0;
    if(execute_CsrPlugin_csr_768) begin
      _zz_CsrPlugin_csrMapping_readDataInit_2[12 : 11] = CsrPlugin_mstatus_MPP;
      _zz_CsrPlugin_csrMapping_readDataInit_2[7 : 7] = CsrPlugin_mstatus_MPIE;
      _zz_CsrPlugin_csrMapping_readDataInit_2[3 : 3] = CsrPlugin_mstatus_MIE;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_3 = 32'h0;
    if(execute_CsrPlugin_csr_836) begin
      _zz_CsrPlugin_csrMapping_readDataInit_3[11 : 11] = CsrPlugin_mip_MEIP;
      _zz_CsrPlugin_csrMapping_readDataInit_3[7 : 7] = CsrPlugin_mip_MTIP;
      _zz_CsrPlugin_csrMapping_readDataInit_3[3 : 3] = CsrPlugin_mip_MSIP;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_4 = 32'h0;
    if(execute_CsrPlugin_csr_772) begin
      _zz_CsrPlugin_csrMapping_readDataInit_4[11 : 11] = CsrPlugin_mie_MEIE;
      _zz_CsrPlugin_csrMapping_readDataInit_4[7 : 7] = CsrPlugin_mie_MTIE;
      _zz_CsrPlugin_csrMapping_readDataInit_4[3 : 3] = CsrPlugin_mie_MSIE;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_5 = 32'h0;
    if(execute_CsrPlugin_csr_833) begin
      _zz_CsrPlugin_csrMapping_readDataInit_5[31 : 0] = CsrPlugin_mepc;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_6 = 32'h0;
    if(execute_CsrPlugin_csr_834) begin
      _zz_CsrPlugin_csrMapping_readDataInit_6[31 : 31] = CsrPlugin_mcause_interrupt;
      _zz_CsrPlugin_csrMapping_readDataInit_6[3 : 0] = CsrPlugin_mcause_exceptionCode;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_7 = 32'h0;
    if(execute_CsrPlugin_csr_835) begin
      _zz_CsrPlugin_csrMapping_readDataInit_7[31 : 0] = CsrPlugin_mtval;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_8 = 32'h0;
    if(execute_CsrPlugin_csr_3008) begin
      _zz_CsrPlugin_csrMapping_readDataInit_8[31 : 0] = _zz_CsrPlugin_csrMapping_readDataInit;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_9 = 32'h0;
    if(execute_CsrPlugin_csr_4032) begin
      _zz_CsrPlugin_csrMapping_readDataInit_9[31 : 0] = _zz_CsrPlugin_csrMapping_readDataInit_1;
    end
  end

  assign CsrPlugin_csrMapping_readDataInit = (((_zz_CsrPlugin_csrMapping_readDataInit_2 | _zz_CsrPlugin_csrMapping_readDataInit_3) | (_zz_CsrPlugin_csrMapping_readDataInit_4 | _zz_CsrPlugin_csrMapping_readDataInit_5)) | ((_zz_CsrPlugin_csrMapping_readDataInit_6 | _zz_CsrPlugin_csrMapping_readDataInit_7) | (_zz_CsrPlugin_csrMapping_readDataInit_8 | _zz_CsrPlugin_csrMapping_readDataInit_9)));
  assign when_CsrPlugin_l1297 = (CsrPlugin_privilege < execute_CsrPlugin_csrAddress[9 : 8]);
  assign when_CsrPlugin_l1302 = ((! execute_arbitration_isValid) || (! execute_IS_CSR));
  assign iBusWishbone_ADR = {_zz_iBusWishbone_ADR_1,_zz_iBusWishbone_ADR};
  assign iBusWishbone_CTI = ((_zz_iBusWishbone_ADR == 3'b111) ? 3'b111 : 3'b010);
  assign iBusWishbone_BTE = 2'b00;
  assign iBusWishbone_SEL = 4'b1111;
  assign iBusWishbone_WE = 1'b0;
  assign iBusWishbone_DAT_MOSI = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  always @(*) begin
    iBusWishbone_CYC = 1'b0;
    if(when_InstructionCache_l239) begin
      iBusWishbone_CYC = 1'b1;
    end
  end

  always @(*) begin
    iBusWishbone_STB = 1'b0;
    if(when_InstructionCache_l239) begin
      iBusWishbone_STB = 1'b1;
    end
  end

  assign when_InstructionCache_l239 = (iBus_cmd_valid || (_zz_iBusWishbone_ADR != 3'b000));
  assign iBus_cmd_ready = (iBus_cmd_valid && iBusWishbone_ACK);
  assign iBus_rsp_valid = _zz_iBus_rsp_valid;
  assign iBus_rsp_payload_data = iBusWishbone_DAT_MISO_regNext;
  assign iBus_rsp_payload_error = 1'b0;
  assign dBus_cmd_halfPipe_fire = (dBus_cmd_halfPipe_valid && dBus_cmd_halfPipe_ready);
  assign dBus_cmd_ready = (! dBus_cmd_rValid);
  assign dBus_cmd_halfPipe_valid = dBus_cmd_rValid;
  assign dBus_cmd_halfPipe_payload_wr = dBus_cmd_rData_wr;
  assign dBus_cmd_halfPipe_payload_address = dBus_cmd_rData_address;
  assign dBus_cmd_halfPipe_payload_data = dBus_cmd_rData_data;
  assign dBus_cmd_halfPipe_payload_size = dBus_cmd_rData_size;
  assign dBusWishbone_ADR = (dBus_cmd_halfPipe_payload_address >>> 2);
  assign dBusWishbone_CTI = 3'b000;
  assign dBusWishbone_BTE = 2'b00;
  always @(*) begin
    case(dBus_cmd_halfPipe_payload_size)
      2'b00 : begin
        _zz_dBusWishbone_SEL = 4'b0001;
      end
      2'b01 : begin
        _zz_dBusWishbone_SEL = 4'b0011;
      end
      default : begin
        _zz_dBusWishbone_SEL = 4'b1111;
      end
    endcase
  end

  always @(*) begin
    dBusWishbone_SEL = (_zz_dBusWishbone_SEL <<< dBus_cmd_halfPipe_payload_address[1 : 0]);
    if(when_DBusSimplePlugin_l189) begin
      dBusWishbone_SEL = 4'b1111;
    end
  end

  assign when_DBusSimplePlugin_l189 = (! dBus_cmd_halfPipe_payload_wr);
  assign dBusWishbone_WE = dBus_cmd_halfPipe_payload_wr;
  assign dBusWishbone_DAT_MOSI = dBus_cmd_halfPipe_payload_data;
  assign dBus_cmd_halfPipe_ready = (dBus_cmd_halfPipe_valid && dBusWishbone_ACK);
  assign dBusWishbone_CYC = dBus_cmd_halfPipe_valid;
  assign dBusWishbone_STB = dBus_cmd_halfPipe_valid;
  assign dBus_rsp_ready = ((dBus_cmd_halfPipe_valid && (! dBusWishbone_WE)) && dBusWishbone_ACK);
  assign dBus_rsp_data = dBusWishbone_DAT_MISO;
  assign dBus_rsp_error = 1'b0;
  always @(posedge clk) begin
    if(reset) begin
      IBusCachedPlugin_fetchPc_pcReg <= externalResetVector;
      IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      IBusCachedPlugin_fetchPc_booted <= 1'b0;
      IBusCachedPlugin_fetchPc_inc <= 1'b0;
      _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= 1'b0;
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      IBusCachedPlugin_rspCounter <= _zz_IBusCachedPlugin_rspCounter;
      IBusCachedPlugin_rspCounter <= 32'h0;
      _zz_2 <= 1'b1;
      execute_LightShifterPlugin_isActive <= 1'b0;
      HazardSimplePlugin_writeBackBuffer_valid <= 1'b0;
      CsrPlugin_mstatus_MIE <= 1'b0;
      CsrPlugin_mstatus_MPIE <= 1'b0;
      CsrPlugin_mstatus_MPP <= 2'b11;
      CsrPlugin_mie_MEIE <= 1'b0;
      CsrPlugin_mie_MTIE <= 1'b0;
      CsrPlugin_mie_MSIE <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      CsrPlugin_interrupt_valid <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      CsrPlugin_hadException <= 1'b0;
      execute_CsrPlugin_wfiWake <= 1'b0;
      _zz_CsrPlugin_csrMapping_readDataInit <= 32'h0;
      execute_arbitration_isValid <= 1'b0;
      memory_arbitration_isValid <= 1'b0;
      writeBack_arbitration_isValid <= 1'b0;
      switch_Fetcher_l362 <= 3'b000;
      _zz_iBusWishbone_ADR <= 3'b000;
      _zz_iBus_rsp_valid <= 1'b0;
      dBus_cmd_rValid <= 1'b0;
    end else begin
      if(IBusCachedPlugin_fetchPc_correction) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b1;
      end
      if(IBusCachedPlugin_fetchPc_output_fire) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      end
      IBusCachedPlugin_fetchPc_booted <= 1'b1;
      if(when_Fetcher_l131) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_output_fire_1) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b1;
      end
      if(when_Fetcher_l131_1) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(when_Fetcher_l158) begin
        IBusCachedPlugin_fetchPc_pcReg <= IBusCachedPlugin_fetchPc_pc;
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= 1'b0;
      end
      if(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= (IBusCachedPlugin_iBusRsp_stages_0_output_valid && (! 1'b0));
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      end
      if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= (IBusCachedPlugin_iBusRsp_stages_1_output_valid && (! IBusCachedPlugin_iBusRsp_flush));
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      end
      if(when_Fetcher_l329) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b1;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      end
      if(when_Fetcher_l329_1) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= IBusCachedPlugin_injector_nextPcCalc_valids_0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      end
      if(when_Fetcher_l329_2) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= IBusCachedPlugin_injector_nextPcCalc_valids_1;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      end
      if(when_Fetcher_l329_3) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= IBusCachedPlugin_injector_nextPcCalc_valids_2;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      end
      if(when_Fetcher_l329_4) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= IBusCachedPlugin_injector_nextPcCalc_valids_3;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      end
      if(iBus_rsp_valid) begin
        IBusCachedPlugin_rspCounter <= (IBusCachedPlugin_rspCounter + 32'h00000001);
      end
      
        


          if(!(! (((dBus_rsp_ready && memory_MEMORY_ENABLE) && memory_arbitration_isValid) && memory_arbitration_isStuck))) begin
            $display("FAILURE DBusSimplePlugin doesn't allow memory stage stall when read happend");
            $finish;
          end
        
      
      
        


          if(!(! (((writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE) && (! writeBack_MEMORY_STORE)) && writeBack_arbitration_isStuck))) begin
            $display("FAILURE DBusSimplePlugin doesn't allow writeback stage stall when read happend");
            $finish;
          end
        
      
      _zz_2 <= 1'b0;
      if(when_ShiftPlugins_l169) begin
        if(when_ShiftPlugins_l175) begin
          execute_LightShifterPlugin_isActive <= 1'b1;
          if(execute_LightShifterPlugin_done) begin
            execute_LightShifterPlugin_isActive <= 1'b0;
          end
        end
      end
      if(execute_arbitration_removeIt) begin
        execute_LightShifterPlugin_isActive <= 1'b0;
      end
      HazardSimplePlugin_writeBackBuffer_valid <= HazardSimplePlugin_writeBackWrites_valid;
      if(when_CsrPlugin_l909) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
      end
      if(when_CsrPlugin_l909_1) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= (CsrPlugin_exceptionPortCtrl_exceptionValids_decode && (! decode_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
      end
      if(when_CsrPlugin_l909_2) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= (CsrPlugin_exceptionPortCtrl_exceptionValids_execute && (! execute_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
      end
      if(when_CsrPlugin_l909_3) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= (CsrPlugin_exceptionPortCtrl_exceptionValids_memory && (! memory_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      end
      CsrPlugin_interrupt_valid <= 1'b0;
      if(when_CsrPlugin_l946) begin
        if(when_CsrPlugin_l952) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l952_1) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l952_2) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
      end
      if(CsrPlugin_pipelineLiberator_active) begin
        if(when_CsrPlugin_l980) begin
          CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b1;
        end
        if(when_CsrPlugin_l980_1) begin
          CsrPlugin_pipelineLiberator_pcValids_1 <= CsrPlugin_pipelineLiberator_pcValids_0;
        end
        if(when_CsrPlugin_l980_2) begin
          CsrPlugin_pipelineLiberator_pcValids_2 <= CsrPlugin_pipelineLiberator_pcValids_1;
        end
      end
      if(when_CsrPlugin_l985) begin
        CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      end
      if(CsrPlugin_interruptJump) begin
        CsrPlugin_interrupt_valid <= 1'b0;
      end
      CsrPlugin_hadException <= CsrPlugin_exception;
      if(when_CsrPlugin_l1019) begin
        case(CsrPlugin_targetPrivilege)
          2'b11 : begin
            CsrPlugin_mstatus_MIE <= 1'b0;
            CsrPlugin_mstatus_MPIE <= CsrPlugin_mstatus_MIE;
            CsrPlugin_mstatus_MPP <= CsrPlugin_privilege;
          end
          default : begin
          end
        endcase
      end
      if(when_CsrPlugin_l1064) begin
        case(switch_CsrPlugin_l1068)
          2'b11 : begin
            CsrPlugin_mstatus_MPP <= 2'b00;
            CsrPlugin_mstatus_MIE <= CsrPlugin_mstatus_MPIE;
            CsrPlugin_mstatus_MPIE <= 1'b1;
          end
          default : begin
          end
        endcase
      end
      execute_CsrPlugin_wfiWake <= (({_zz_when_CsrPlugin_l952_2,{_zz_when_CsrPlugin_l952_1,_zz_when_CsrPlugin_l952}} != 3'b000) || CsrPlugin_thirdPartyWake);
      if(when_Pipeline_l151) begin
        execute_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154) begin
        execute_arbitration_isValid <= decode_arbitration_isValid;
      end
      if(when_Pipeline_l151_1) begin
        memory_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_1) begin
        memory_arbitration_isValid <= execute_arbitration_isValid;
      end
      if(when_Pipeline_l151_2) begin
        writeBack_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_2) begin
        writeBack_arbitration_isValid <= memory_arbitration_isValid;
      end
      case(switch_Fetcher_l362)
        3'b000 : begin
          if(IBusCachedPlugin_injectionPort_valid) begin
            switch_Fetcher_l362 <= 3'b001;
          end
        end
        3'b001 : begin
          switch_Fetcher_l362 <= 3'b010;
        end
        3'b010 : begin
          switch_Fetcher_l362 <= 3'b011;
        end
        3'b011 : begin
          if(when_Fetcher_l378) begin
            switch_Fetcher_l362 <= 3'b100;
          end
        end
        3'b100 : begin
          switch_Fetcher_l362 <= 3'b000;
        end
        default : begin
        end
      endcase
      if(execute_CsrPlugin_csr_768) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mstatus_MPP <= CsrPlugin_csrMapping_writeDataSignal[12 : 11];
          CsrPlugin_mstatus_MPIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mstatus_MIE <= CsrPlugin_csrMapping_writeDataSignal[3];
        end
      end
      if(execute_CsrPlugin_csr_772) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mie_MEIE <= CsrPlugin_csrMapping_writeDataSignal[11];
          CsrPlugin_mie_MTIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mie_MSIE <= CsrPlugin_csrMapping_writeDataSignal[3];
        end
      end
      if(execute_CsrPlugin_csr_3008) begin
        if(execute_CsrPlugin_writeEnable) begin
          _zz_CsrPlugin_csrMapping_readDataInit <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
        end
      end
      if(when_InstructionCache_l239) begin
        if(iBusWishbone_ACK) begin
          _zz_iBusWishbone_ADR <= (_zz_iBusWishbone_ADR + 3'b001);
        end
      end
      _zz_iBus_rsp_valid <= (iBusWishbone_CYC && iBusWishbone_ACK);
      if(dBus_cmd_valid) begin
        dBus_cmd_rValid <= 1'b1;
      end
      if(dBus_cmd_halfPipe_fire) begin
        dBus_cmd_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload <= IBusCachedPlugin_iBusRsp_stages_1_output_payload;
    end
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_s1_tightlyCoupledHit <= IBusCachedPlugin_s0_tightlyCoupledHit;
    end
    if(IBusCachedPlugin_iBusRsp_stages_2_input_ready) begin
      IBusCachedPlugin_s2_tightlyCoupledHit <= IBusCachedPlugin_s1_tightlyCoupledHit;
    end
    if(when_ShiftPlugins_l169) begin
      if(when_ShiftPlugins_l175) begin
        execute_LightShifterPlugin_amplitudeReg <= (execute_LightShifterPlugin_amplitude - 5'h01);
      end
    end
    HazardSimplePlugin_writeBackBuffer_payload_address <= HazardSimplePlugin_writeBackWrites_payload_address;
    HazardSimplePlugin_writeBackBuffer_payload_data <= HazardSimplePlugin_writeBackWrites_payload_data;
    CsrPlugin_mip_MEIP <= externalInterrupt;
    CsrPlugin_mip_MTIP <= timerInterrupt;
    CsrPlugin_mip_MSIP <= softwareInterrupt;
    CsrPlugin_mcycle <= (CsrPlugin_mcycle + 64'h0000000000000001);
    if(writeBack_arbitration_isFiring) begin
      CsrPlugin_minstret <= (CsrPlugin_minstret + 64'h0000000000000001);
    end
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_code : decodeExceptionPort_payload_code);
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_badAddr : decodeExceptionPort_payload_badAddr);
    end
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= CsrPlugin_selfException_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= CsrPlugin_selfException_payload_badAddr;
    end
    if(_zz_when_1) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3 ? DBusSimplePlugin_memoryExceptionPort_payload_code : BranchPlugin_branchExceptionPort_payload_code);
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_3 ? DBusSimplePlugin_memoryExceptionPort_payload_badAddr : BranchPlugin_branchExceptionPort_payload_badAddr);
    end
    if(when_CsrPlugin_l946) begin
      if(when_CsrPlugin_l952) begin
        CsrPlugin_interrupt_code <= 4'b0111;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l952_1) begin
        CsrPlugin_interrupt_code <= 4'b0011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l952_2) begin
        CsrPlugin_interrupt_code <= 4'b1011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
    end
    if(when_CsrPlugin_l1019) begin
      case(CsrPlugin_targetPrivilege)
        2'b11 : begin
          CsrPlugin_mcause_interrupt <= (! CsrPlugin_hadException);
          CsrPlugin_mcause_exceptionCode <= CsrPlugin_trapCause;
          CsrPlugin_mepc <= writeBack_PC;
          if(CsrPlugin_hadException) begin
            CsrPlugin_mtval <= CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
          end
        end
        default : begin
        end
      endcase
    end
    externalInterruptArray_regNext <= externalInterruptArray;
    if(when_Pipeline_l124) begin
      decode_to_execute_PC <= decode_PC;
    end
    if(when_Pipeline_l124_1) begin
      execute_to_memory_PC <= _zz_execute_SRC2;
    end
    if(when_Pipeline_l124_2) begin
      memory_to_writeBack_PC <= memory_PC;
    end
    if(when_Pipeline_l124_3) begin
      decode_to_execute_INSTRUCTION <= decode_INSTRUCTION;
    end
    if(when_Pipeline_l124_4) begin
      execute_to_memory_INSTRUCTION <= execute_INSTRUCTION;
    end
    if(when_Pipeline_l124_5) begin
      memory_to_writeBack_INSTRUCTION <= memory_INSTRUCTION;
    end
    if(when_Pipeline_l124_6) begin
      decode_to_execute_FORMAL_PC_NEXT <= decode_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_7) begin
      execute_to_memory_FORMAL_PC_NEXT <= execute_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_8) begin
      memory_to_writeBack_FORMAL_PC_NEXT <= _zz_memory_to_writeBack_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_9) begin
      decode_to_execute_SRC1_CTRL <= _zz_decode_to_execute_SRC1_CTRL;
    end
    if(when_Pipeline_l124_10) begin
      decode_to_execute_SRC_USE_SUB_LESS <= decode_SRC_USE_SUB_LESS;
    end
    if(when_Pipeline_l124_11) begin
      decode_to_execute_MEMORY_ENABLE <= decode_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_12) begin
      execute_to_memory_MEMORY_ENABLE <= execute_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_13) begin
      memory_to_writeBack_MEMORY_ENABLE <= memory_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_14) begin
      decode_to_execute_ALU_CTRL <= _zz_decode_to_execute_ALU_CTRL;
    end
    if(when_Pipeline_l124_15) begin
      decode_to_execute_SRC2_CTRL <= _zz_decode_to_execute_SRC2_CTRL;
    end
    if(when_Pipeline_l124_16) begin
      decode_to_execute_REGFILE_WRITE_VALID <= decode_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_17) begin
      execute_to_memory_REGFILE_WRITE_VALID <= execute_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_18) begin
      memory_to_writeBack_REGFILE_WRITE_VALID <= memory_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_19) begin
      decode_to_execute_BYPASSABLE_EXECUTE_STAGE <= decode_BYPASSABLE_EXECUTE_STAGE;
    end
    if(when_Pipeline_l124_20) begin
      decode_to_execute_BYPASSABLE_MEMORY_STAGE <= decode_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_21) begin
      execute_to_memory_BYPASSABLE_MEMORY_STAGE <= execute_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_22) begin
      decode_to_execute_MEMORY_STORE <= decode_MEMORY_STORE;
    end
    if(when_Pipeline_l124_23) begin
      execute_to_memory_MEMORY_STORE <= execute_MEMORY_STORE;
    end
    if(when_Pipeline_l124_24) begin
      memory_to_writeBack_MEMORY_STORE <= memory_MEMORY_STORE;
    end
    if(when_Pipeline_l124_25) begin
      decode_to_execute_SRC_LESS_UNSIGNED <= decode_SRC_LESS_UNSIGNED;
    end
    if(when_Pipeline_l124_26) begin
      decode_to_execute_ALU_BITWISE_CTRL <= _zz_decode_to_execute_ALU_BITWISE_CTRL;
    end
    if(when_Pipeline_l124_27) begin
      decode_to_execute_SHIFT_CTRL <= _zz_decode_to_execute_SHIFT_CTRL;
    end
    if(when_Pipeline_l124_28) begin
      decode_to_execute_BRANCH_CTRL <= _zz_decode_to_execute_BRANCH_CTRL;
    end
    if(when_Pipeline_l124_29) begin
      decode_to_execute_IS_CSR <= decode_IS_CSR;
    end
    if(when_Pipeline_l124_30) begin
      decode_to_execute_ENV_CTRL <= _zz_decode_to_execute_ENV_CTRL;
    end
    if(when_Pipeline_l124_31) begin
      execute_to_memory_ENV_CTRL <= _zz_execute_to_memory_ENV_CTRL;
    end
    if(when_Pipeline_l124_32) begin
      memory_to_writeBack_ENV_CTRL <= _zz_memory_to_writeBack_ENV_CTRL;
    end
    if(when_Pipeline_l124_33) begin
      decode_to_execute_RS1 <= decode_RS1;
    end
    if(when_Pipeline_l124_34) begin
      decode_to_execute_RS2 <= decode_RS2;
    end
    if(when_Pipeline_l124_35) begin
      decode_to_execute_SRC2_FORCE_ZERO <= decode_SRC2_FORCE_ZERO;
    end
    if(when_Pipeline_l124_36) begin
      decode_to_execute_CSR_WRITE_OPCODE <= decode_CSR_WRITE_OPCODE;
    end
    if(when_Pipeline_l124_37) begin
      decode_to_execute_CSR_READ_OPCODE <= decode_CSR_READ_OPCODE;
    end
    if(when_Pipeline_l124_38) begin
      decode_to_execute_DO_EBREAK <= decode_DO_EBREAK;
    end
    if(when_Pipeline_l124_39) begin
      execute_to_memory_ALIGNEMENT_FAULT <= execute_ALIGNEMENT_FAULT;
    end
    if(when_Pipeline_l124_40) begin
      execute_to_memory_MEMORY_ADDRESS_LOW <= execute_MEMORY_ADDRESS_LOW;
    end
    if(when_Pipeline_l124_41) begin
      memory_to_writeBack_MEMORY_ADDRESS_LOW <= memory_MEMORY_ADDRESS_LOW;
    end
    if(when_Pipeline_l124_42) begin
      execute_to_memory_REGFILE_WRITE_DATA <= _zz_execute_to_memory_REGFILE_WRITE_DATA;
    end
    if(when_Pipeline_l124_43) begin
      memory_to_writeBack_REGFILE_WRITE_DATA <= memory_REGFILE_WRITE_DATA;
    end
    if(when_Pipeline_l124_44) begin
      execute_to_memory_BRANCH_DO <= execute_BRANCH_DO;
    end
    if(when_Pipeline_l124_45) begin
      execute_to_memory_BRANCH_CALC <= execute_BRANCH_CALC;
    end
    if(when_Pipeline_l124_46) begin
      memory_to_writeBack_MEMORY_READ_DATA <= memory_MEMORY_READ_DATA;
    end
    if(when_CsrPlugin_l1264) begin
      execute_CsrPlugin_csr_768 <= (decode_INSTRUCTION[31 : 20] == 12'h300);
    end
    if(when_CsrPlugin_l1264_1) begin
      execute_CsrPlugin_csr_836 <= (decode_INSTRUCTION[31 : 20] == 12'h344);
    end
    if(when_CsrPlugin_l1264_2) begin
      execute_CsrPlugin_csr_772 <= (decode_INSTRUCTION[31 : 20] == 12'h304);
    end
    if(when_CsrPlugin_l1264_3) begin
      execute_CsrPlugin_csr_773 <= (decode_INSTRUCTION[31 : 20] == 12'h305);
    end
    if(when_CsrPlugin_l1264_4) begin
      execute_CsrPlugin_csr_833 <= (decode_INSTRUCTION[31 : 20] == 12'h341);
    end
    if(when_CsrPlugin_l1264_5) begin
      execute_CsrPlugin_csr_834 <= (decode_INSTRUCTION[31 : 20] == 12'h342);
    end
    if(when_CsrPlugin_l1264_6) begin
      execute_CsrPlugin_csr_835 <= (decode_INSTRUCTION[31 : 20] == 12'h343);
    end
    if(when_CsrPlugin_l1264_7) begin
      execute_CsrPlugin_csr_3008 <= (decode_INSTRUCTION[31 : 20] == 12'hbc0);
    end
    if(when_CsrPlugin_l1264_8) begin
      execute_CsrPlugin_csr_4032 <= (decode_INSTRUCTION[31 : 20] == 12'hfc0);
    end
    if(execute_CsrPlugin_csr_836) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mip_MSIP <= CsrPlugin_csrMapping_writeDataSignal[3];
      end
    end
    if(execute_CsrPlugin_csr_773) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mtvec_base <= CsrPlugin_csrMapping_writeDataSignal[31 : 2];
        CsrPlugin_mtvec_mode <= CsrPlugin_csrMapping_writeDataSignal[1 : 0];
      end
    end
    if(execute_CsrPlugin_csr_833) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mepc <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    iBusWishbone_DAT_MISO_regNext <= iBusWishbone_DAT_MISO;
    if(dBus_cmd_ready) begin
      dBus_cmd_rData_wr <= dBus_cmd_payload_wr;
      dBus_cmd_rData_address <= dBus_cmd_payload_address;
      dBus_cmd_rData_data <= dBus_cmd_payload_data;
      dBus_cmd_rData_size <= dBus_cmd_payload_size;
    end
  end

  always @(posedge clk) begin
    DebugPlugin_firstCycle <= 1'b0;
    if(debug_bus_cmd_ready) begin
      DebugPlugin_firstCycle <= 1'b1;
    end
    DebugPlugin_secondCycle <= DebugPlugin_firstCycle;
    DebugPlugin_isPipBusy <= (({writeBack_arbitration_isValid,{memory_arbitration_isValid,{execute_arbitration_isValid,decode_arbitration_isValid}}} != 4'b0000) || IBusCachedPlugin_incomingInstruction);
    if(writeBack_arbitration_isValid) begin
      DebugPlugin_busReadDataReg <= _zz_lastStageRegFileWrite_payload_data;
    end
    _zz_when_DebugPlugin_l244 <= debug_bus_cmd_payload_address[2];
    if(when_DebugPlugin_l284) begin
      DebugPlugin_busReadDataReg <= execute_PC;
    end
    DebugPlugin_resetIt_regNext <= DebugPlugin_resetIt;
  end

  always @(posedge clk) begin
    if(debugReset) begin
      DebugPlugin_resetIt <= 1'b0;
      DebugPlugin_haltIt <= 1'b0;
      DebugPlugin_stepIt <= 1'b0;
      DebugPlugin_godmode <= 1'b0;
      DebugPlugin_haltedByBreak <= 1'b0;
      DebugPlugin_debugUsed <= 1'b0;
      DebugPlugin_disableEbreak <= 1'b0;
    end else begin
      if(when_DebugPlugin_l225) begin
        DebugPlugin_godmode <= 1'b1;
      end
      if(debug_bus_cmd_valid) begin
        DebugPlugin_debugUsed <= 1'b1;
      end
      if(debug_bus_cmd_valid) begin
        case(switch_DebugPlugin_l256)
          6'h0 : begin
            if(debug_bus_cmd_payload_wr) begin
              DebugPlugin_stepIt <= debug_bus_cmd_payload_data[4];
              if(when_DebugPlugin_l260) begin
                DebugPlugin_resetIt <= 1'b1;
              end
              if(when_DebugPlugin_l260_1) begin
                DebugPlugin_resetIt <= 1'b0;
              end
              if(when_DebugPlugin_l261) begin
                DebugPlugin_haltIt <= 1'b1;
              end
              if(when_DebugPlugin_l261_1) begin
                DebugPlugin_haltIt <= 1'b0;
              end
              if(when_DebugPlugin_l262) begin
                DebugPlugin_haltedByBreak <= 1'b0;
              end
              if(when_DebugPlugin_l263) begin
                DebugPlugin_godmode <= 1'b0;
              end
              if(when_DebugPlugin_l264) begin
                DebugPlugin_disableEbreak <= 1'b1;
              end
              if(when_DebugPlugin_l264_1) begin
                DebugPlugin_disableEbreak <= 1'b0;
              end
            end
          end
          default : begin
          end
        endcase
      end
      if(when_DebugPlugin_l284) begin
        if(when_DebugPlugin_l287) begin
          DebugPlugin_haltIt <= 1'b1;
          DebugPlugin_haltedByBreak <= 1'b1;
        end
      end
      if(when_DebugPlugin_l300) begin
        if(decode_arbitration_isValid) begin
          DebugPlugin_haltIt <= 1'b1;
        end
      end
    end
  end


endmodule

module InstructionCache (
  input               io_flush,
  input               io_cpu_prefetch_isValid,
  output reg          io_cpu_prefetch_haltIt,
  input      [31:0]   io_cpu_prefetch_pc,
  input               io_cpu_fetch_isValid,
  input               io_cpu_fetch_isStuck,
  input               io_cpu_fetch_isRemoved,
  input      [31:0]   io_cpu_fetch_pc,
  output     [31:0]   io_cpu_fetch_data,
  input      [31:0]   io_cpu_fetch_mmuRsp_physicalAddress,
  input               io_cpu_fetch_mmuRsp_isIoAccess,
  input               io_cpu_fetch_mmuRsp_isPaging,
  input               io_cpu_fetch_mmuRsp_allowRead,
  input               io_cpu_fetch_mmuRsp_allowWrite,
  input               io_cpu_fetch_mmuRsp_allowExecute,
  input               io_cpu_fetch_mmuRsp_exception,
  input               io_cpu_fetch_mmuRsp_refilling,
  input               io_cpu_fetch_mmuRsp_bypassTranslation,
  output     [31:0]   io_cpu_fetch_physicalAddress,
  input               io_cpu_decode_isValid,
  input               io_cpu_decode_isStuck,
  input      [31:0]   io_cpu_decode_pc,
  output     [31:0]   io_cpu_decode_physicalAddress,
  output     [31:0]   io_cpu_decode_data,
  output              io_cpu_decode_cacheMiss,
  output              io_cpu_decode_error,
  output              io_cpu_decode_mmuRefilling,
  output              io_cpu_decode_mmuException,
  input               io_cpu_decode_isUser,
  input               io_cpu_fill_valid,
  input      [31:0]   io_cpu_fill_payload,
  output              io_mem_cmd_valid,
  input               io_mem_cmd_ready,
  output     [31:0]   io_mem_cmd_payload_address,
  output     [2:0]    io_mem_cmd_payload_size,
  input               io_mem_rsp_valid,
  input      [31:0]   io_mem_rsp_payload_data,
  input               io_mem_rsp_payload_error,
  input      [2:0]    _zz_when_Fetcher_l398,
  input      [31:0]   _zz_io_cpu_fetch_data_regNextWhen,
  input               clk,
  input               reset
);
  reg        [31:0]   _zz_banks_0_port1;
  reg        [27:0]   _zz_ways_0_tags_port1;
  wire       [27:0]   _zz_ways_0_tags_port;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 lineLoader_fire;
  reg                 lineLoader_valid;
  (* keep , syn_keep *) reg        [31:0]   lineLoader_address /* synthesis syn_keep = 1 */ ;
  reg                 lineLoader_hadError;
  reg                 lineLoader_flushPending;
  reg        [1:0]    lineLoader_flushCounter;
  wire                when_InstructionCache_l338;
  reg                 _zz_when_InstructionCache_l342;
  wire                when_InstructionCache_l342;
  wire                when_InstructionCache_l351;
  reg                 lineLoader_cmdSent;
  wire                io_mem_cmd_fire;
  wire                when_Utils_l357;
  reg                 lineLoader_wayToAllocate_willIncrement;
  wire                lineLoader_wayToAllocate_willClear;
  wire                lineLoader_wayToAllocate_willOverflowIfInc;
  wire                lineLoader_wayToAllocate_willOverflow;
  (* keep , syn_keep *) reg        [2:0]    lineLoader_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                lineLoader_write_tag_0_valid;
  wire       [0:0]    lineLoader_write_tag_0_payload_address;
  wire                lineLoader_write_tag_0_payload_data_valid;
  wire                lineLoader_write_tag_0_payload_data_error;
  wire       [25:0]   lineLoader_write_tag_0_payload_data_address;
  wire                lineLoader_write_data_0_valid;
  wire       [3:0]    lineLoader_write_data_0_payload_address;
  wire       [31:0]   lineLoader_write_data_0_payload_data;
  wire                when_InstructionCache_l401;
  wire       [3:0]    _zz_fetchStage_read_banksValue_0_dataMem;
  wire                _zz_fetchStage_read_banksValue_0_dataMem_1;
  wire       [31:0]   fetchStage_read_banksValue_0_dataMem;
  wire       [31:0]   fetchStage_read_banksValue_0_data;
  wire       [0:0]    _zz_fetchStage_read_waysValues_0_tag_valid;
  wire                _zz_fetchStage_read_waysValues_0_tag_valid_1;
  wire                fetchStage_read_waysValues_0_tag_valid;
  wire                fetchStage_read_waysValues_0_tag_error;
  wire       [25:0]   fetchStage_read_waysValues_0_tag_address;
  wire       [27:0]   _zz_fetchStage_read_waysValues_0_tag_valid_2;
  wire                fetchStage_hit_hits_0;
  wire                fetchStage_hit_valid;
  wire                fetchStage_hit_error;
  wire       [31:0]   fetchStage_hit_data;
  wire       [31:0]   fetchStage_hit_word;
  wire                when_InstructionCache_l435;
  reg        [31:0]   io_cpu_fetch_data_regNextWhen;
  wire                when_InstructionCache_l459;
  reg        [31:0]   decodeStage_mmuRsp_physicalAddress;
  reg                 decodeStage_mmuRsp_isIoAccess;
  reg                 decodeStage_mmuRsp_isPaging;
  reg                 decodeStage_mmuRsp_allowRead;
  reg                 decodeStage_mmuRsp_allowWrite;
  reg                 decodeStage_mmuRsp_allowExecute;
  reg                 decodeStage_mmuRsp_exception;
  reg                 decodeStage_mmuRsp_refilling;
  reg                 decodeStage_mmuRsp_bypassTranslation;
  wire                when_InstructionCache_l459_1;
  reg                 decodeStage_hit_valid;
  wire                when_InstructionCache_l459_2;
  reg                 decodeStage_hit_error;
  wire                when_Fetcher_l398;
  (* ram_style = "block" *) reg [31:0] banks_0 [0:15];
  (* ram_style = "block" *) reg [27:0] ways_0_tags [0:1];

  assign _zz_ways_0_tags_port = {lineLoader_write_tag_0_payload_data_address,{lineLoader_write_tag_0_payload_data_error,lineLoader_write_tag_0_payload_data_valid}};
  always @(posedge clk) begin
    if(_zz_1) begin
      banks_0[lineLoader_write_data_0_payload_address] <= lineLoader_write_data_0_payload_data;
    end
  end

  always @(posedge clk) begin
    if(_zz_fetchStage_read_banksValue_0_dataMem_1) begin
      _zz_banks_0_port1 <= banks_0[_zz_fetchStage_read_banksValue_0_dataMem];
    end
  end

  always @(posedge clk) begin
    if(_zz_2) begin
      ways_0_tags[lineLoader_write_tag_0_payload_address] <= _zz_ways_0_tags_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_fetchStage_read_waysValues_0_tag_valid_1) begin
      _zz_ways_0_tags_port1 <= ways_0_tags[_zz_fetchStage_read_waysValues_0_tag_valid];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(lineLoader_write_data_0_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(lineLoader_write_tag_0_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    lineLoader_fire = 1'b0;
    if(io_mem_rsp_valid) begin
      if(when_InstructionCache_l401) begin
        lineLoader_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    io_cpu_prefetch_haltIt = (lineLoader_valid || lineLoader_flushPending);
    if(when_InstructionCache_l338) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
    if(when_InstructionCache_l342) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
    if(io_flush) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
  end

  assign when_InstructionCache_l338 = (! lineLoader_flushCounter[1]);
  assign when_InstructionCache_l342 = (! _zz_when_InstructionCache_l342);
  assign when_InstructionCache_l351 = (lineLoader_flushPending && (! (lineLoader_valid || io_cpu_fetch_isValid)));
  assign io_mem_cmd_fire = (io_mem_cmd_valid && io_mem_cmd_ready);
  assign io_mem_cmd_valid = (lineLoader_valid && (! lineLoader_cmdSent));
  assign io_mem_cmd_payload_address = {lineLoader_address[31 : 5],5'h0};
  assign io_mem_cmd_payload_size = 3'b101;
  assign when_Utils_l357 = (! lineLoader_valid);
  always @(*) begin
    lineLoader_wayToAllocate_willIncrement = 1'b0;
    if(when_Utils_l357) begin
      lineLoader_wayToAllocate_willIncrement = 1'b1;
    end
  end

  assign lineLoader_wayToAllocate_willClear = 1'b0;
  assign lineLoader_wayToAllocate_willOverflowIfInc = 1'b1;
  assign lineLoader_wayToAllocate_willOverflow = (lineLoader_wayToAllocate_willOverflowIfInc && lineLoader_wayToAllocate_willIncrement);
  assign lineLoader_write_tag_0_valid = ((1'b1 && lineLoader_fire) || (! lineLoader_flushCounter[1]));
  assign lineLoader_write_tag_0_payload_address = (lineLoader_flushCounter[1] ? lineLoader_address[5 : 5] : lineLoader_flushCounter[0 : 0]);
  assign lineLoader_write_tag_0_payload_data_valid = lineLoader_flushCounter[1];
  assign lineLoader_write_tag_0_payload_data_error = (lineLoader_hadError || io_mem_rsp_payload_error);
  assign lineLoader_write_tag_0_payload_data_address = lineLoader_address[31 : 6];
  assign lineLoader_write_data_0_valid = (io_mem_rsp_valid && 1'b1);
  assign lineLoader_write_data_0_payload_address = {lineLoader_address[5 : 5],lineLoader_wordIndex};
  assign lineLoader_write_data_0_payload_data = io_mem_rsp_payload_data;
  assign when_InstructionCache_l401 = (lineLoader_wordIndex == 3'b111);
  assign _zz_fetchStage_read_banksValue_0_dataMem = io_cpu_prefetch_pc[5 : 2];
  assign _zz_fetchStage_read_banksValue_0_dataMem_1 = (! io_cpu_fetch_isStuck);
  assign fetchStage_read_banksValue_0_dataMem = _zz_banks_0_port1;
  assign fetchStage_read_banksValue_0_data = fetchStage_read_banksValue_0_dataMem[31 : 0];
  assign _zz_fetchStage_read_waysValues_0_tag_valid = io_cpu_prefetch_pc[5 : 5];
  assign _zz_fetchStage_read_waysValues_0_tag_valid_1 = (! io_cpu_fetch_isStuck);
  assign _zz_fetchStage_read_waysValues_0_tag_valid_2 = _zz_ways_0_tags_port1;
  assign fetchStage_read_waysValues_0_tag_valid = _zz_fetchStage_read_waysValues_0_tag_valid_2[0];
  assign fetchStage_read_waysValues_0_tag_error = _zz_fetchStage_read_waysValues_0_tag_valid_2[1];
  assign fetchStage_read_waysValues_0_tag_address = _zz_fetchStage_read_waysValues_0_tag_valid_2[27 : 2];
  assign fetchStage_hit_hits_0 = (fetchStage_read_waysValues_0_tag_valid && (fetchStage_read_waysValues_0_tag_address == io_cpu_fetch_mmuRsp_physicalAddress[31 : 6]));
  assign fetchStage_hit_valid = (fetchStage_hit_hits_0 != 1'b0);
  assign fetchStage_hit_error = fetchStage_read_waysValues_0_tag_error;
  assign fetchStage_hit_data = fetchStage_read_banksValue_0_data;
  assign fetchStage_hit_word = fetchStage_hit_data;
  assign io_cpu_fetch_data = fetchStage_hit_word;
  assign when_InstructionCache_l435 = (! io_cpu_decode_isStuck);
  assign io_cpu_decode_data = io_cpu_fetch_data_regNextWhen;
  assign io_cpu_fetch_physicalAddress = io_cpu_fetch_mmuRsp_physicalAddress;
  assign when_InstructionCache_l459 = (! io_cpu_decode_isStuck);
  assign when_InstructionCache_l459_1 = (! io_cpu_decode_isStuck);
  assign when_InstructionCache_l459_2 = (! io_cpu_decode_isStuck);
  assign io_cpu_decode_cacheMiss = (! decodeStage_hit_valid);
  assign io_cpu_decode_error = (decodeStage_hit_error || ((! decodeStage_mmuRsp_isPaging) && (decodeStage_mmuRsp_exception || (! decodeStage_mmuRsp_allowExecute))));
  assign io_cpu_decode_mmuRefilling = decodeStage_mmuRsp_refilling;
  assign io_cpu_decode_mmuException = (((! decodeStage_mmuRsp_refilling) && decodeStage_mmuRsp_isPaging) && (decodeStage_mmuRsp_exception || (! decodeStage_mmuRsp_allowExecute)));
  assign io_cpu_decode_physicalAddress = decodeStage_mmuRsp_physicalAddress;
  assign when_Fetcher_l398 = (_zz_when_Fetcher_l398 != 3'b000);
  always @(posedge clk) begin
    if(reset) begin
      lineLoader_valid <= 1'b0;
      lineLoader_hadError <= 1'b0;
      lineLoader_flushPending <= 1'b1;
      lineLoader_cmdSent <= 1'b0;
      lineLoader_wordIndex <= 3'b000;
    end else begin
      if(lineLoader_fire) begin
        lineLoader_valid <= 1'b0;
      end
      if(lineLoader_fire) begin
        lineLoader_hadError <= 1'b0;
      end
      if(io_cpu_fill_valid) begin
        lineLoader_valid <= 1'b1;
      end
      if(io_flush) begin
        lineLoader_flushPending <= 1'b1;
      end
      if(when_InstructionCache_l351) begin
        lineLoader_flushPending <= 1'b0;
      end
      if(io_mem_cmd_fire) begin
        lineLoader_cmdSent <= 1'b1;
      end
      if(lineLoader_fire) begin
        lineLoader_cmdSent <= 1'b0;
      end
      if(io_mem_rsp_valid) begin
        lineLoader_wordIndex <= (lineLoader_wordIndex + 3'b001);
        if(io_mem_rsp_payload_error) begin
          lineLoader_hadError <= 1'b1;
        end
      end
    end
  end

  always @(posedge clk) begin
    if(io_cpu_fill_valid) begin
      lineLoader_address <= io_cpu_fill_payload;
    end
    if(when_InstructionCache_l338) begin
      lineLoader_flushCounter <= (lineLoader_flushCounter + 2'b01);
    end
    _zz_when_InstructionCache_l342 <= lineLoader_flushCounter[1];
    if(when_InstructionCache_l351) begin
      lineLoader_flushCounter <= 2'b00;
    end
    if(when_InstructionCache_l435) begin
      io_cpu_fetch_data_regNextWhen <= io_cpu_fetch_data;
    end
    if(when_InstructionCache_l459) begin
      decodeStage_mmuRsp_physicalAddress <= io_cpu_fetch_mmuRsp_physicalAddress;
      decodeStage_mmuRsp_isIoAccess <= io_cpu_fetch_mmuRsp_isIoAccess;
      decodeStage_mmuRsp_isPaging <= io_cpu_fetch_mmuRsp_isPaging;
      decodeStage_mmuRsp_allowRead <= io_cpu_fetch_mmuRsp_allowRead;
      decodeStage_mmuRsp_allowWrite <= io_cpu_fetch_mmuRsp_allowWrite;
      decodeStage_mmuRsp_allowExecute <= io_cpu_fetch_mmuRsp_allowExecute;
      decodeStage_mmuRsp_exception <= io_cpu_fetch_mmuRsp_exception;
      decodeStage_mmuRsp_refilling <= io_cpu_fetch_mmuRsp_refilling;
      decodeStage_mmuRsp_bypassTranslation <= io_cpu_fetch_mmuRsp_bypassTranslation;
    end
    if(when_InstructionCache_l459_1) begin
      decodeStage_hit_valid <= fetchStage_hit_valid;
    end
    if(when_InstructionCache_l459_2) begin
      decodeStage_hit_error <= fetchStage_hit_error;
    end
    if(when_Fetcher_l398) begin
      io_cpu_fetch_data_regNextWhen <= _zz_io_cpu_fetch_data_regNextWhen;
    end
  end


endmodule
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// `default_nettype none
 
	













	













	

































































































































































// `default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

















































 // __GLOBAL_DEFINE_H
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none


// User GPIO initial configuration parameters


// Useful GPIO mode values.  These match the names used in defs.h.















// The power-on configuration for GPIO 0 to 4 is fixed and cannot be
// modified (allowing the SPI and debug to always be accessible unless
// overridden by a flash program).

// The values below can be any of the standard types defined above,
// or they can be any 13-bit value if the user wants a non-standard
// startup state for the GPIO.  By default, every GPIO from 5 to 37
// is set to power up as an input controlled by the management SoC.
// Users may want to redefine these so that the user project powers
// up in a state that can be used immediately without depending on
// the management SoC to run a startup program to configure the GPIOs.











// Configurations of GPIO 14 to 24 are used on caravel but not caravan.


























 // __USER_DEFINES_H
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// `default_nettype none

/* Define the array of GPIO pads.  Note that the analog project support
 * version of caravel (caravan) defines fewer GPIO and replaces them
 * with analog in the chip_io_alt module.  Because the pad signalling
 * remains the same, `MPRJ_IO_PADS does not change, so a local parameter
 * is made that can be made smaller than `MPRJ_IO_PADS to accommodate
 * the analog pads.
 */

module mprj_io #(
    parameter AREA1PADS = 19,
    parameter TOTAL_PADS = (19 + 19)
) (
    inout vddio,
    inout vssio,
    inout vdda,
    inout vssa,
    inout vccd,
    inout vssd,

    inout vdda1,
    inout vdda2,
    inout vssa1,
    inout vssa2,

    input vddio_q,
    input vssio_q,
    input analog_a,
    input analog_b,
    input porb_h,
    input [TOTAL_PADS-1:0] vccd_conb,
    inout [TOTAL_PADS-1:0] io,
    input [TOTAL_PADS-1:0] io_out,
    input [TOTAL_PADS-1:0] oeb,
    input [TOTAL_PADS-1:0] enh,
    input [TOTAL_PADS-1:0] inp_dis,
    input [TOTAL_PADS-1:0] ib_mode_sel,
    input [TOTAL_PADS-1:0] vtrip_sel,
    input [TOTAL_PADS-1:0] slow_sel,
    input [TOTAL_PADS-1:0] holdover,
    input [TOTAL_PADS-1:0] analog_en,
    input [TOTAL_PADS-1:0] analog_sel,
    input [TOTAL_PADS-1:0] analog_pol,
    input [TOTAL_PADS*3-1:0] dm,
    output [TOTAL_PADS-1:0] io_in,
    output [TOTAL_PADS-1:0] io_in_3v3,
    inout [TOTAL_PADS-10:0] analog_io,
    inout [TOTAL_PADS-10:0] analog_noesd_io
);

    wire [TOTAL_PADS-1:0] loop0_io;	// Internal loopback to 3.3V domain ground
    wire [TOTAL_PADS-1:0] loop1_io;	// Internal loopback to 3.3V domain power
    wire [6:0] no_connect_1a, no_connect_1b;
    wire [1:0] no_connect_2a, no_connect_2b;

    sky130_ef_io__gpiov2_pad_wrapped  area1_io_pad [AREA1PADS - 1:0] (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
	    .PAD(io[AREA1PADS - 1:0]),
	
	    .OUT(io_out[AREA1PADS - 1:0]),
	    .OE_N(oeb[AREA1PADS - 1:0]),
	    .HLD_H_N(loop1_io[AREA1PADS - 1:0]),
	    .ENABLE_H(enh[AREA1PADS - 1:0]),
	    .ENABLE_INP_H(loop0_io[AREA1PADS - 1:0]),
	    .ENABLE_VDDA_H(porb_h),
	    .ENABLE_VSWITCH_H(loop0_io[AREA1PADS - 1:0]),
	    .ENABLE_VDDIO(vccd_conb[AREA1PADS - 1:0]),
	    .INP_DIS(inp_dis[AREA1PADS - 1:0]),
	    .IB_MODE_SEL(ib_mode_sel[AREA1PADS - 1:0]),
	    .VTRIP_SEL(vtrip_sel[AREA1PADS - 1:0]),
	    .SLOW(slow_sel[AREA1PADS - 1:0]),
	    .HLD_OVR(holdover[AREA1PADS - 1:0]),
	    .ANALOG_EN(analog_en[AREA1PADS - 1:0]),
	    .ANALOG_SEL(analog_sel[AREA1PADS - 1:0]),
	    .ANALOG_POL(analog_pol[AREA1PADS - 1:0]),
	    .DM(dm[AREA1PADS*3 - 1:0]),
	    .PAD_A_NOESD_H({analog_noesd_io[AREA1PADS - 8:0], no_connect_1a}),
	    .PAD_A_ESD_0_H({analog_io[AREA1PADS - 8:0], no_connect_1b}),
	    .PAD_A_ESD_1_H(),
	    .IN(io_in[AREA1PADS - 1:0]),
	    .IN_H(io_in_3v3[AREA1PADS - 1:0]),
	    .TIE_HI_ESD(loop1_io[AREA1PADS - 1:0]),
	    .TIE_LO_ESD(loop0_io[AREA1PADS - 1:0])
    );

    sky130_ef_io__gpiov2_pad_wrapped area2_io_pad [TOTAL_PADS - AREA1PADS - 1:0] (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
	    .PAD(io[TOTAL_PADS - 1:AREA1PADS]),
	
	    .OUT(io_out[TOTAL_PADS - 1:AREA1PADS]),
	    .OE_N(oeb[TOTAL_PADS - 1:AREA1PADS]),
	    .HLD_H_N(loop1_io[TOTAL_PADS - 1:AREA1PADS]),
	    .ENABLE_H(enh[TOTAL_PADS - 1:AREA1PADS]),
	    .ENABLE_INP_H(loop0_io[TOTAL_PADS - 1:AREA1PADS]),
	    .ENABLE_VDDA_H(porb_h),
	    .ENABLE_VSWITCH_H(loop0_io[TOTAL_PADS - 1:AREA1PADS]),
	    .ENABLE_VDDIO(vccd_conb[TOTAL_PADS - 1:AREA1PADS]),
	    .INP_DIS(inp_dis[TOTAL_PADS - 1:AREA1PADS]),
	    .IB_MODE_SEL(ib_mode_sel[TOTAL_PADS - 1:AREA1PADS]),
	    .VTRIP_SEL(vtrip_sel[TOTAL_PADS - 1:AREA1PADS]),
	    .SLOW(slow_sel[TOTAL_PADS - 1:AREA1PADS]),
	    .HLD_OVR(holdover[TOTAL_PADS - 1:AREA1PADS]),
	    .ANALOG_EN(analog_en[TOTAL_PADS - 1:AREA1PADS]),
	    .ANALOG_SEL(analog_sel[TOTAL_PADS - 1:AREA1PADS]),
	    .ANALOG_POL(analog_pol[TOTAL_PADS - 1:AREA1PADS]),
	    .DM(dm[TOTAL_PADS*3 - 1:AREA1PADS*3]),
	    .PAD_A_NOESD_H({no_connect_2a, analog_noesd_io[TOTAL_PADS - 10:AREA1PADS - 7]}),
	    .PAD_A_ESD_0_H({no_connect_2b, analog_io[TOTAL_PADS - 10:AREA1PADS - 7]}),
	    .PAD_A_ESD_1_H(),
	    .IN(io_in[TOTAL_PADS - 1:AREA1PADS]),
	    .IN_H(io_in_3v3[TOTAL_PADS - 1:AREA1PADS]),
	    .TIE_HI_ESD(loop1_io[TOTAL_PADS - 1:AREA1PADS]),
	    .TIE_LO_ESD(loop0_io[TOTAL_PADS - 1:AREA1PADS])
    );

endmodule
// `default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
`timescale 1 ns / 1 ps

module simple_por(

    inout vdd3v3,
    inout vdd1v8,
    inout vss3v3,
    inout vss1v8,

    output porb_h,
    output porb_l,
    output por_l
);

    wire mid;
    reg inode;

    // This is a behavioral model!  Actual circuit is a resitor dumping
    // current (slowly) from vdd3v3 onto a capacitor, and this fed into
    // two schmitt triggers for strong hysteresis/glitch tolerance.

    initial begin
	inode <= 1'b0; 
    end 

    // Emulate current source on capacitor as a 500ns delay either up or
    // down.  Note that this is sped way up for verilog simulation;  the
    // actual circuit is set to a 15ms delay.

    always @(posedge vdd3v3) begin
	#500 inode <= 1'b1;
    end
    always @(negedge vdd3v3) begin
	#500 inode <= 1'b0;
    end

    // Instantiate two shmitt trigger buffers in series

    sky130_fd_sc_hvl__schmittbuf_1 hystbuf1 (

	.VPWR(vdd3v3),
	.VGND(vss3v3),
	.VPB(vdd3v3),
	.VNB(vss3v3),

	.A(inode),
	.X(mid)
    );

    sky130_fd_sc_hvl__schmittbuf_1 hystbuf2 (

	.VPWR(vdd3v3),
	.VGND(vss3v3),
	.VPB(vdd3v3),
	.VNB(vss3v3),

	.A(mid),
	.X(porb_h)
    );

    sky130_fd_sc_hvl__lsbufhv2lv_1 porb_level (

	.VPWR(vdd3v3),
	.VPB(vdd3v3),
	.LVPWR(vdd1v8),
	.VNB(vss3v3),
	.VGND(vss3v3),

	.A(porb_h),
	.X(porb_l)
    );

    // since this is behavioral anyway, but this should be
    // replaced by a proper inverter
    assign por_l = ~porb_l;
endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
// (True) digital PLL
//
// Output goes to a trimmable ring oscillator (see documentation).
// Ring oscillator should be trimmable to above and below maximum
// ranges of the input.
//
// Input "osc" comes from a fixed clock source (e.g., crystal oscillator
// output).
//
// Input "div" is the target number of clock cycles per oscillator cycle.
// e.g., if div == 8 then this is an 8X PLL.
//
// Clock "clock" is the PLL output being trimmed.
// (NOTE:  To be done:  Pass-through enable)
//
// Algorithm:
//
// 1) Trim is done by thermometer code.  Reset to the highest value
//    in case the fastest rate clock is too fast for the logic.
//
// 2) Count the number of contiguous 1s and 0s in "osc"
//    periods of the master clock.  If the count maxes out, it does
//    not roll over.
//
// 3) Add the two counts together.
//
// 4) If the sum is less than div, then the clock is too slow, so
//    decrease the trim code.  If the sum is greater than div, the
//    clock is too fast, so increase the trim code.  If the sum
//    is equal to div, the the trim code does not change.
//

module digital_pll_controller(reset, clock, osc, div, trim);
    input reset;
    input clock;
    input osc;
    input [4:0] div;
    output [25:0] trim;		// Use ring_osc2x13, with 26 trim bits

    wire [25:0] trim;
    reg [2:0] oscbuf;
    reg [2:0] prep;

    reg [4:0] count0;
    reg [4:0] count1;
    reg [6:0] tval;	// Includes 2 bits fractional
    wire [4:0] tint;	// Integer part of the above

    wire [5:0] sum;

    assign sum = count0 + count1;
 
    // Integer to thermometer code (maybe there's an algorithmic way?)
    assign tint = tval[6:2];
                                     // |<--second-->|<-- first-->|
    assign trim = (tint == 5'd0)  ? 26'b0000000000000_0000000000000 :
          (tint == 5'd1)  ? 26'b0000000000000_0000000000001 :
          (tint == 5'd2)  ? 26'b0000000000000_0000001000001 :
          (tint == 5'd3)  ? 26'b0000000000000_0010001000001 :
          (tint == 5'd4)  ? 26'b0000000000000_0010001001001 :
          (tint == 5'd5)  ? 26'b0000000000000_0010101001001 :
          (tint == 5'd6)  ? 26'b0000000000000_1010101001001 :
          (tint == 5'd7)  ? 26'b0000000000000_1010101101001 :
          (tint == 5'd8)  ? 26'b0000000000000_1010101101101 :
          (tint == 5'd9)  ? 26'b0000000000000_1011101101101 :
          (tint == 5'd10) ? 26'b0000000000000_1011101111101 :
          (tint == 5'd11) ? 26'b0000000000000_1111101111101 :
          (tint == 5'd12) ? 26'b0000000000000_1111101111111 :
          (tint == 5'd13) ? 26'b0000000000000_1111111111111 :
          (tint == 5'd14) ? 26'b0000000000001_1111111111111 :
          (tint == 5'd15) ? 26'b0000001000001_1111111111111 :
          (tint == 5'd16) ? 26'b0010001000001_1111111111111 :
          (tint == 5'd17) ? 26'b0010001001001_1111111111111 :
          (tint == 5'd18) ? 26'b0010101001001_1111111111111 :
          (tint == 5'd19) ? 26'b1010101001001_1111111111111 :
          (tint == 5'd20) ? 26'b1010101101001_1111111111111 :
          (tint == 5'd21) ? 26'b1010101101101_1111111111111 :
          (tint == 5'd22) ? 26'b1011101101101_1111111111111 :
          (tint == 5'd23) ? 26'b1011101111101_1111111111111 :
          (tint == 5'd24) ? 26'b1111101111101_1111111111111 :
          (tint == 5'd25) ? 26'b1111101111111_1111111111111 :
                    26'b1111111111111_1111111111111;
   
    always @(posedge clock or posedge reset) begin
    if (reset == 1'b1) begin
        tval <= 7'd0;	// Note:  trim[0] must be zero for startup to work.
        oscbuf <= 3'd0;
        prep <= 3'd0;
        count0 <= 5'd0;
        count1 <= 5'd0;

    end else begin
        oscbuf <= {oscbuf[1:0], osc};

        if (oscbuf[2] != oscbuf[1]) begin
        count1 <= count0;
        count0 <= 5'b00001;
        prep <= {prep[1:0], 1'b1};

        if (prep == 3'b111) begin
            if (sum > div) begin
		if (tval < 127) begin
            	    tval <= tval + 1;
		end
            end else if (sum < div) begin
		if (tval > 0) begin
            	    tval <= tval - 1;
		end
            end
        end
        end else begin
        if (count0 != 5'b11111) begin
                count0 <= count0 + 1;
        end
        end
    end
    end

endmodule	// digital_pll_controller
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
// Tunable ring oscillator---synthesizable (physical) version.
//
// NOTE:  This netlist cannot be simulated correctly due to lack
// of accurate timing in the digital cell verilog models.

module delay_stage(in, trim, out);
    input in;
    input [1:0] trim;
    output out;

    wire d0, d1, d2, ts;

    sky130_fd_sc_hd__clkbuf_2 delaybuf0 (
	.A(in),
	.X(ts)
    );

    sky130_fd_sc_hd__clkbuf_1 delaybuf1 (
	.A(ts),
	.X(d0)
    );

    sky130_fd_sc_hd__einvp_2 delayen1 (
	.A(d0),
	.TE(trim[1]),
	.Z(d1)
    );

    sky130_fd_sc_hd__einvn_4 delayenb1 (
	.A(ts),
	.TE_B(trim[1]),
	.Z(d1)
    );

    sky130_fd_sc_hd__clkinv_1 delayint0 (
	.A(d1),
	.Y(d2)
    );

    sky130_fd_sc_hd__einvp_2 delayen0 (
	.A(d2),
	.TE(trim[0]),
	.Z(out)
    );

    sky130_fd_sc_hd__einvn_8 delayenb0 (
	.A(ts),
	.TE_B(trim[0]),
	.Z(out)
    );

endmodule

module start_stage(in, trim, reset, out);
    input in;
    input [1:0] trim;
    input reset;
    output out;

    wire d0, d1, d2, ctrl0, one;

    sky130_fd_sc_hd__clkbuf_1 delaybuf0 (
	.A(in),
	.X(d0)
    );

    sky130_fd_sc_hd__einvp_2 delayen1 (
	.A(d0),
	.TE(trim[1]),
	.Z(d1)
    );

    sky130_fd_sc_hd__einvn_4 delayenb1 (
	.A(in),
	.TE_B(trim[1]),
	.Z(d1)
    );

    sky130_fd_sc_hd__clkinv_1 delayint0 (
	.A(d1),
	.Y(d2)
    );

    sky130_fd_sc_hd__einvp_2 delayen0 (
	.A(d2),
	.TE(trim[0]),
	.Z(out)
    );

    sky130_fd_sc_hd__einvn_8 delayenb0 (
	.A(in),
	.TE_B(ctrl0),
	.Z(out)
    );

    sky130_fd_sc_hd__einvp_1 reseten0 (
	.A(one),
	.TE(reset),
	.Z(out)
    );

    sky130_fd_sc_hd__or2_2 ctrlen0 (
	.A(reset),
	.B(trim[0]),
	.X(ctrl0)
    );

    sky130_fd_sc_hd__conb_1 const1 (
	.HI(one),
	.LO()
    );

endmodule

// Ring oscillator with 13 stages, each with two trim bits delay
// (see above).  Trim is not binary:  For trim[1:0], lower bit
// trim[0] is primary trim and must be applied first;  upper
// bit trim[1] is secondary trim and should only be applied
// after the primary trim is applied, or it has no effect.
//
// Total effective number of inverter stages in this oscillator
// ranges from 13 at trim 0 to 65 at trim 24.  The intention is
// to cover a range greater than 2x so that the midrange can be
// reached over all PVT conditions.
//
// Frequency of this ring oscillator under SPICE simulations at
// nominal PVT is maximum 214 MHz (trim 0), minimum 90 MHz (trim 24).

module ring_osc2x13(reset, trim, clockp);
    input reset;
    input [25:0] trim;
    output[1:0] clockp;

	// i.e., behavioral model below

    reg [1:0] clockp;
    reg hiclock;
    integer i;
    real delay;
    wire [5:0] bcount;

    assign bcount = trim[0] + trim[1] + trim[2]
		+ trim[3] + trim[4] + trim[5] + trim[6] + trim[7]
		+ trim[8] + trim[9] + trim[10] + trim[11] + trim[12]
		+ trim[13] + trim[14] + trim[15] + trim[16] + trim[17]
		+ trim[18] + trim[19] + trim[20] + trim[21] + trim[22]
		+ trim[23] + trim[24] + trim[25];

    initial begin
	hiclock <= 1'b0;
	delay = 3.0;
    end

    // Fastest operation is 214 MHz = 4.67ns
    // Delay per trim is 0.02385
    // Run "hiclock" at 2x this rate, then use positive and negative
    // edges to derive the 0 and 90 degree phase clocks.

    always #delay begin
	hiclock <= (hiclock === 1'b0);
    end

    always @(trim) begin
    	// Implement trim as a variable delay, one delay per trim bit
	delay = 1.168 + 0.012 * $itor(bcount);
    end

    always @(posedge hiclock or posedge reset) begin
	if (reset == 1'b1) begin
	    clockp[0] <= 1'b0;
	end else begin
	    clockp[0] <= (clockp[0] === 1'b0);
	end
    end

    always @(negedge hiclock or posedge reset) begin
	if (reset == 1'b1) begin
	    clockp[1] <= 1'b0;
	end else begin
	    clockp[1] <= (clockp[1] === 1'b0);
	end
    end
















































 // !FUNCTIONAL

endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Integer-N clock divider */
`default_nettype none
 
module clock_div #(
    parameter SIZE = 3		// Number of bits for the divider value
) (
    in, out, N, resetb
);
    input in;			// input clock
    input [SIZE-1:0] N;		// the number to be divided by
    input resetb;		// asynchronous reset (sense negative)
    output out;			// divided output clock
 
    wire out_odd;		// output of odd divider
    wire out_even;		// output of even divider
    wire not_zero;		// signal to find divide by 0 case
    wire enable_even;		// enable of even divider
    wire enable_odd;		// enable of odd divider

    reg [SIZE-1:0] syncN;	// N synchronized to output clock
    reg [SIZE-1:0] syncNp;	// N synchronized to output clock
 
    assign not_zero = | syncN[SIZE-1:1];
 
    assign out = (out_odd & syncN[0] & not_zero) | (out_even & !syncN[0]);
    assign enable_odd = syncN[0] & not_zero;
    assign enable_even = !syncN[0];

    // Divider value synchronization (double-synchronized to avoid metastability)
    always @(posedge out or negedge resetb) begin
	if (resetb == 1'b0) begin
	    syncN <= 3'b010;	// Default to divide-by-2 on system reset
	    syncNp <= 3'b010;	// Default to divide-by-2 on system reset
	end else begin
	    syncNp <= N;
	    syncN <= syncNp;
	end
    end
 
    // Even divider
    even even_0(in, out_even, syncN, resetb, not_zero, enable_even);
    // Odd divider
    odd odd_0(in, out_odd, syncN, resetb, enable_odd);
 
endmodule // clock_div
 
/* Odd divider */

module odd #(
    parameter SIZE = 3
) (
    clk, out, N, resetb, enable
);
    input clk;			// slow clock
    output out;			// fast output clock
    input [SIZE-1:0] N;		// division factor
    input resetb;		// synchronous reset
    input enable;		// odd enable
 
    reg [SIZE-1:0] counter;	// these 2 counters are used
    reg [SIZE-1:0] counter2;	// to non-overlapping signals
    reg out_counter;		// positive edge triggered counter
    reg out_counter2;		// negative edge triggered counter
    reg rst_pulse;		// pulse generated when vector N changes
    reg [SIZE-1:0] old_N;	// gets set to old N when N is changed
    wire not_zero;		// if !not_zero, we devide by 1
 
    // xor to generate 50% duty, half-period waves of final output
    assign out = out_counter2 ^ out_counter;

    // positive edge counter/divider
    always @(posedge clk or negedge resetb) begin
	if (resetb == 1'b0) begin
	    counter <= 3'b010;
	    out_counter <= 1;
	end else if (rst_pulse) begin
	    counter <= N;
	    out_counter <= 1;
	end else if (enable) begin
	    if (counter == 1) begin
		counter <= N;
		out_counter <= ~out_counter;
	    end else begin
		counter <= counter - 1'b1;
	    end
	end
    end
 
    reg [SIZE-1:0] initial_begin;	// this is used to offset the negative edge counter
    wire [SIZE:0] interm_3;		// from the positive edge counter in order to
    assign interm_3 = {1'b0, N} + 2'b11;	// guarantee 50% duty cycle.

    localparam [SIZE:0] interm_init = {1'b0,3'b010} + 2'b11;

    // Counter driven by negative edge of clock.

    always @(negedge clk or negedge resetb) begin
	if (resetb == 1'b0) begin
	    // reset the counter at system reset
	    counter2 <= 3'b010;
	    initial_begin <= interm_init[SIZE:1];
	    out_counter2 <= 1;
	end else if (rst_pulse) begin
	    // reset the counter at change of N.
	    counter2 <= N;
	    initial_begin <= interm_3[SIZE:1];
	    out_counter2 <= 1;
	end else if ((initial_begin <= 1) && enable) begin

	    // Do normal logic after odd calibration.
	    // This is the same as the even counter.
	    if (counter2 == 1) begin
		counter2 <= N;
		out_counter2 <= ~out_counter2;
	    end else begin
		counter2 <= counter2 - 1'b1;
	    end
	end else if (enable) begin
	    initial_begin <= initial_begin - 1'b1;
	end
    end
 
    //
    // reset pulse generator:
    //               __    __    __    __    _
    // clk:       __/  \__/  \__/  \__/  \__/
    //            _ __________________________
    // N:         _X__________________________
    //               _____
    // rst_pulse: __/     \___________________
    //
    // This block generates an internal reset for the odd divider in the
    // form of a single pulse signal when the odd divider is enabled.

    always @(posedge clk or negedge resetb) begin
	if (resetb == 1'b0) begin
	    rst_pulse <= 0;
	end else if (enable) begin
	    if (N != old_N) begin
		// pulse when reset changes
		rst_pulse <= 1;
	    end else begin
		rst_pulse <= 0;
	    end
	end
    end
 
    always @(posedge clk) begin
	// always save the old N value to guarante reset from
	// an even-to-odd transition.
	old_N <= N;
    end	
 
endmodule // odd

/* Even divider */

module even #(
    parameter SIZE = 3
) (
    clk, out, N, resetb, not_zero, enable
);
    input clk;		// fast input clock
    output out;		// slower divided clock
    input [SIZE-1:0] N;	// divide by factor 'N'
    input resetb;	// asynchronous reset
    input not_zero;	// if !not_zero divide by 1
    input enable;	// enable the even divider
 
    reg [SIZE-1:0] counter;
    reg out_counter;
    wire [SIZE-1:0] div_2;
 
    // if N=0 just output the clock, otherwise, divide it.
    assign out = (clk & !not_zero) | (out_counter & not_zero);
    assign div_2 = {1'b0, N[SIZE-1:1]};
 
    // simple flip-flop even divider
    always @(posedge clk or negedge resetb) begin
	if (resetb == 1'b0) begin
	    counter <= 1;
	    out_counter <= 1;

	end else if (enable) begin
	    // only use switching power if enabled
	    if (counter == 1) begin
		// divide after counter has reached bottom
		// of interval 'N' which will be value '1'
		counter <= div_2;
		out_counter <= ~out_counter;
	    end else begin
		// decrement the counter and wait
		counter <= counter-1;	// to start next transition.
	    end
	end
    end
 
endmodule //even
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

//-----------------------------------------------------------
// SPI controller for Caravel
//-----------------------------------------------------------
// housekeeping_spi.v
//------------------------------------------------------
// General purpose SPI module for the Caravel chip
//------------------------------------------------------
// Written by Tim Edwards
// efabless, inc., September 28, 2020
//------------------------------------------------
// This file is distributed free and open source
//------------------------------------------------

// SCK ---   Clock input
// SDI ---   Data  input
// SDO ---   Data  output
// CSB ---   Chip  select (sense negative)
// idata --- Data from chip to transmit out, in 8 bits
// odata --- Input data to chip, in 8 bits
// addr  --- Decoded address to upstream circuits
// rdstb --- Read strobe, tells upstream circuit that data will be latched.
// wrstb --- Write strobe, tells upstream circuit to latch odata.

// Data format (general purpose):
// 8 bit format
// 1st byte:   Command word (see below)
// 2nd byte:   Address word (register 0 to 255)
// 3rd byte:   Data word    (value 0 to 255)

// Command format:
// 00000000  No operation
// 10000000  Write until CSB raised
// 01000000  Read  until CSB raised
// 11000000  Simultaneous read/write until CSB raised
// 11000100  Pass-through read/write to management area flash SPI until CSB raised
// 11000010  Pass-through read/write to user area flash SPI until CSB raised
// wrnnn000  Read/write as above, for nnn = 1 to 7 bytes, then terminate

// Lower three bits are reserved for future use.
// All serial bytes are read and written msb first.

// Fixed control and status registers

// Address 0 is reserved and contains flags for SPI mode.  This is
// currently undefined and is always value 0.
// Address 1 is reserved and contains manufacturer ID low 8 bits.
// Address 2 is reserved and contains manufacturer ID high 4 bits.
// Address 3 is reserved and contains product ID (8 bits).
// Addresses 4 to 7 are reserved and contain the mask ID (32 bits).
// Addresses 8 to 255 are available for general purpose use.







module housekeeping_spi(reset, SCK, SDI, CSB, SDO,
	sdoenb, idata, odata, oaddr, rdstb, wrstb,
	pass_thru_mgmt, pass_thru_mgmt_delay,
	pass_thru_user, pass_thru_user_delay,
	pass_thru_mgmt_reset, pass_thru_user_reset);

    input reset;
    input SCK;
    input SDI;
    input CSB;
    output SDO;
    output sdoenb;
    input [7:0] idata;
    output [7:0] odata;
    output [7:0] oaddr;
    output rdstb;
    output wrstb; 
    output pass_thru_mgmt;
    output pass_thru_mgmt_delay;
    output pass_thru_user;
    output pass_thru_user_delay;
    output pass_thru_mgmt_reset;
    output pass_thru_user_reset;

    reg  [7:0]  addr;
    reg		wrstb;
    reg		rdstb;
    reg		sdoenb;
    reg  [2:0]  state;
    reg  [2:0]  count;
    reg		writemode;
    reg		readmode;
    reg  [2:0]	fixed;
    wire [7:0]  odata;
    reg  [6:0]  predata;
    wire [7:0]  oaddr;
    reg  [7:0]  ldata;
    reg		pass_thru_mgmt;
    reg		pass_thru_mgmt_delay;
    reg		pre_pass_thru_mgmt;
    reg		pass_thru_user;
    reg		pass_thru_user_delay;
    reg		pre_pass_thru_user;
    wire	csb_reset;

    assign odata = {predata, SDI};
    assign oaddr = (state == 3'b001) ? {addr[6:0], SDI} : addr;
    assign SDO = ldata[7];
    assign csb_reset = CSB | reset;
    assign pass_thru_mgmt_reset = pass_thru_mgmt_delay | pre_pass_thru_mgmt;
    assign pass_thru_user_reset = pass_thru_user_delay | pre_pass_thru_user;

    // Readback data is captured on the falling edge of SCK so that
    // it is guaranteed valid at the next rising edge.
    always @(negedge SCK or posedge csb_reset) begin
        if (csb_reset == 1'b1) begin
            wrstb <= 1'b0;
            ldata  <= 8'b00000000;
            sdoenb <= 1'b1;
        end else begin

            // After CSB low, 1st SCK starts command

            if (state == 3'b010) begin
            	if (readmode == 1'b1) begin
                    sdoenb <= 1'b0;
                    if (count == 3'b000) begin
                	ldata <= idata;
                    end else begin
                	ldata <= {ldata[6:0], 1'b0};	// Shift out
                    end
                end else begin
                    sdoenb <= 1'b1;
                end

                // Apply write strobe on SCK negative edge on the next-to-last
                // data bit so that it updates data on the rising edge of SCK
                // on the last data bit.
 
                if (count == 3'b111) begin
                    if (writemode == 1'b1) begin
                        wrstb <= 1'b1;
                    end
                end else begin
                    wrstb <= 1'b0;
                end

	    end else if (state == 3'b101 || state == 3'b100) begin
		wrstb <= 1'b0;
		sdoenb <= 1'b0;
            end else begin
                wrstb <= 1'b0;
                sdoenb <= 1'b1;
            end		// ! state `DATA
        end		// ! csb_reset
    end			// always @ ~SCK

    always @(posedge SCK or posedge csb_reset) begin
        if (csb_reset == 1'b1) begin
            // Default state on reset
            addr <= 8'h00;
	    rdstb <= 1'b0;
            predata <= 7'b0000000;
            state  <= 3'b000;
            count  <= 3'b000;
            readmode <= 1'b0;
            writemode <= 1'b0;
            fixed <= 3'b000;
	    pass_thru_mgmt <= 1'b0;
	    pass_thru_mgmt_delay <= 1'b0;
	    pre_pass_thru_mgmt <= 1'b0;
	    pass_thru_user <= 1'b0;
	    pass_thru_user_delay <= 1'b0;
	    pre_pass_thru_user <= 1'b0;
        end else begin
            // After csb_reset low, 1st SCK starts command
            if (state == 3'b000) begin
		rdstb <= 1'b0;
                count <= count + 1;
        	if (count == 3'b000) begin
	            writemode <= SDI;
	        end else if (count == 3'b001) begin
	            readmode <= SDI;
	        end else if (count < 3'b101) begin
	            fixed <= {fixed[1:0], SDI}; 
	        end else if (count == 3'b101) begin
		    pre_pass_thru_mgmt <= SDI;
	        end else if (count == 3'b110) begin
		    pre_pass_thru_user <= SDI;
		    pass_thru_mgmt_delay <= pre_pass_thru_mgmt;
	        end else if (count == 3'b111) begin
		    pass_thru_user_delay <= pre_pass_thru_user;
		    if (pre_pass_thru_mgmt == 1'b1) begin
			state <= 3'b101;
			pre_pass_thru_mgmt <= 1'b0;
		    end else if (pre_pass_thru_user == 1'b1) begin
			state <= 3'b100;
			pre_pass_thru_user <= 1'b0;
		    end else begin
	                state <= 3'b001;
		    end
	        end
            end else if (state == 3'b001) begin
	        count <= count + 1;
	        addr <= {addr[6:0], SDI};
	        if (count == 3'b111) begin
	            state <= 3'b010;
		    if (readmode == 1'b1) begin
			rdstb <= 1'b1;
		    end
	        end else begin
		    rdstb <= 1'b0;
		end

            end else if (state == 3'b010) begin
	        predata <= {predata[6:0], SDI};
	        count <= count + 1;
	        if (count == 3'b111) begin
	            if (fixed == 3'b001) begin
	                state <= 3'b000;
	            end else if (fixed != 3'b000) begin
	                fixed <= fixed - 1;
	                addr <= addr + 1;	// Auto increment address (fixed)
	            end else begin	
	                addr <= addr + 1;	// Auto increment address (streaming)
	            end
		    if (readmode == 1'b1) begin
			rdstb <= 1'b1;
		    end
	        end else begin
		    rdstb <= 1'b0;
		end
	    end else if (state == 3'b101) begin
		pass_thru_mgmt <= 1'b1;
	    end else if (state == 3'b100) begin
		pass_thru_user <= 1'b1;
            end		// ! state `DATA | `MGMTPASS | `USERPASS
        end		// ! csb_reset 
    end			// always @ SCK

endmodule // housekeeping_spi
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// `default_nettype none

/* Alternative padframe that removes the GPIO from the top row,	*/
/* replacing them with un-overlaid power pads which have a	*/
/* direct connection from pad to core.				*/

/* For convenience, all of the original GPIO signals remain	*/
/* defined in the I/O list, although some are not connected.	*/

/* ANALOG_PADS_1 = Number of GPIO pads in the user 1 section 	*/
/* 		   that are replaced by straight-through analog	*/
/* ANALOG_PADS_2 = Number of GPIO pads in the user 2 section 	*/
/* 		   that are replaced by straight-through analog	*/

module chip_io_alt #(
	parameter ANALOG_PADS_1 = 5,
	parameter ANALOG_PADS_2 = 6
) (
	// Package Pins
	inout  vddio_pad,			// Common padframe/ESD supply
	inout  vddio_pad2,			// Common padframe/ESD supply
	inout  vssio_pad,			// Common padframe/ESD ground
	inout  vssio_pad2,			// Common padframe/ESD ground
	inout  vccd_pad,			// Common 1.8V supply
	inout  vssd_pad,			// Common digital ground
	inout  vdda_pad,			// Management analog 3.3V supply
	inout  vssa_pad,			// Management analog ground
	inout  vdda1_pad,			// User area 1 3.3V supply
	inout  vdda1_pad2,			// User area 1 3.3V supply
	inout  vdda2_pad,			// User area 2 3.3V supply
	inout  vssa1_pad,			// User area 1 analog ground
	inout  vssa1_pad2,			// User area 1 analog ground
	inout  vssa2_pad,			// User area 2 analog ground
	inout  vccd1_pad,			// User area 1 1.8V supply
	inout  vccd2_pad,			// User area 2 1.8V supply
	inout  vssd1_pad,			// User area 1 digital ground
	inout  vssd2_pad,			// User area 2 digital ground

	// Core Side
	inout  vddio,		// Common padframe/ESD supply
	inout  vssio,		// Common padframe/ESD ground
	inout  vccd,		// Common 1.8V supply
	inout  vssd,		// Common digital ground
	inout  vdda,		// Management analog 3.3V supply
	inout  vssa,		// Management analog ground
	inout  vdda1,		// User area 1 3.3V supply
	inout  vdda2,		// User area 2 3.3V supply
	inout  vssa1,		// User area 1 analog ground
	inout  vssa2,		// User area 2 analog ground
	inout  vccd1,		// User area 1 1.8V supply
	inout  vccd2,		// User area 2 1.8V supply
	inout  vssd1,		// User area 1 digital ground
	inout  vssd2,		// User area 2 digital ground

	inout  gpio,
	input  clock,
	input  resetb,
	output flash_csb,
	output flash_clk,
	inout  flash_io0,
	inout  flash_io1,
	// Chip Core Interface
	input  porb_h,
	input  por,
	output resetb_core_h,
	output clock_core,
	input  gpio_out_core,
	output gpio_in_core,
	input  gpio_mode0_core,
	input  gpio_mode1_core,
	input  gpio_outenb_core,
	input  gpio_inenb_core,
	input  flash_csb_core,
	input  flash_clk_core,
	input  flash_csb_oeb_core,
	input  flash_clk_oeb_core,
	input  flash_io0_oeb_core,
	input  flash_io1_oeb_core,
	input  flash_io0_ieb_core,
	input  flash_io1_ieb_core,
	input  flash_io0_do_core,
	input  flash_io1_do_core,
	output flash_io0_di_core,
	output flash_io1_di_core,
	// User project IOs
	// mprj_io is defined for all pads, both digital and analog
	inout [(19 + 19)-1:0] mprj_io,
	// The section below is for the digital pads only.
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_out,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_oeb,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_inp_dis,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_ib_mode_sel,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_vtrip_sel,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_slow_sel,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_holdover,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_analog_en,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_analog_sel,
	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_analog_pol,
	input [((19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2)*3-1:0] mprj_io_dm,
	output [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_in,
	output [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_in_3v3,
 	input [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_one,

	// User project direct access to gpio pad connections for analog
	// "analog" connects to the "esd_0" pin of the GPIO pad, and
	// "analog_noesd" connects to the "noesd" pin of the GPIO pad.

	// User side 1:  Connects to all but the first 7 pads;
	// User side 2:  Connects to all but the last 2 pads
	inout [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-10:0] mprj_gpio_analog,
	inout [(19 + 19)-ANALOG_PADS_1-ANALOG_PADS_2-10:0] mprj_gpio_noesd,

	// Core connections for the analog signals
	inout [ANALOG_PADS_1+ANALOG_PADS_2-1:0] mprj_analog,

	// These are clamp connections for the clamps in the analog cells, if
	// they are used for power supplies.
	// User side 1:  Connects to 
	input [2:0] mprj_clamp_high,
	input [2:0] mprj_clamp_low
);

	wire analog_a, analog_b;
	wire vddio_q, vssio_q;

    // To be considered:  Master hold signal on all user pads (?)
    // For now, set holdh_n to 1 internally (NOTE:  This is in the
    // VDDIO 3.3V domain) and setting enh to porb_h.

    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_enh;

    assign mprj_io_enh = {(19 + 19){porb_h}};

	// Instantiate power and ground pads for management domain
	// 12 pads:  vddio, vssio, vdda, vssa, vccd, vssd
	// One each HV and LV clamp.

	// HV clamps connect between one HV power rail and one ground
	// LV clamps have two clamps connecting between any two LV power
	// rails and grounds, and one back-to-back diode which connects
	// between the first LV clamp ground and any other ground.

    	sky130_ef_io__vddio_hvc_clamped_pad \mgmt_vddio_hvclamp_pad[0]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDIO_PAD(vddio_pad)
    
		);

	// lies in user area 2
    	sky130_ef_io__vddio_hvc_clamped_pad \mgmt_vddio_hvclamp_pad[1]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDIO_PAD(vddio_pad2)

    	);

    	sky130_ef_io__vdda_hvc_clamped_pad mgmt_vdda_hvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDA_PAD(vdda_pad)

	);

    	sky130_ef_io__vccd_lvc_clamped_pad mgmt_vccd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VCCD_PAD(vccd_pad)
    
		);

    	sky130_ef_io__vssio_hvc_clamped_pad \mgmt_vssio_hvclamp_pad[0]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSIO_PAD(vssio_pad)
    
    	);

    	sky130_ef_io__vssio_hvc_clamped_pad \mgmt_vssio_hvclamp_pad[1]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSIO_PAD(vssio_pad2)

    	);

    	sky130_ef_io__vssa_hvc_clamped_pad mgmt_vssa_hvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSA_PAD(vssa_pad)

    	);

    	sky130_ef_io__vssd_lvc_clamped_pad mgmt_vssd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSD_PAD(vssd_pad)

	 	);

	// Instantiate power and ground pads for user 1 domain
	// 8 pads:  vdda, vssa, vccd, vssd;  One each HV and LV clamp.

    	sky130_ef_io__vdda_hvc_clamped_pad \user1_vdda_hvclamp_pad[0] (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDA_PAD(vdda1_pad)

    	);

	    sky130_ef_io__vdda_hvc_clamped_pad \user1_vdda_hvclamp_pad[1] (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDA_PAD(vdda1_pad2)

    	);

    	sky130_ef_io__vccd_lvc_clamped3_pad user1_vccd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		.VCCD1(vccd1),
		.VSSD1(vssd1),

		.VCCD_PAD(vccd1_pad)

    	);

    	sky130_ef_io__vssa_hvc_clamped_pad \user1_vssa_hvclamp_pad[0] (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSA_PAD(vssa1_pad)

    	);

		sky130_ef_io__vssa_hvc_clamped_pad \user1_vssa_hvclamp_pad[1] (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSA_PAD(vssa1_pad2)

    	);

    	sky130_ef_io__vssd_lvc_clamped3_pad user1_vssd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		.VCCD1(vccd1),
		.VSSD1(vssd1),

		.VSSD_PAD(vssd1_pad)

    	);

	// Instantiate power and ground pads for user 2 domain
	// 8 pads:  vdda, vssa, vccd, vssd;  One each HV and LV clamp.

    	sky130_ef_io__vdda_hvc_clamped_pad user2_vdda_hvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDA_PAD(vdda2_pad)

    	);

    	sky130_ef_io__vccd_lvc_clamped3_pad user2_vccd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		.VCCD1(vccd2),
		.VSSD1(vssd2),

		.VCCD_PAD(vccd2_pad)

    	);

    	sky130_ef_io__vssa_hvc_clamped_pad user2_vssa_hvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSA_PAD(vssa2_pad)

    	);

    	sky130_ef_io__vssd_lvc_clamped3_pad user2_vssd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		.VCCD1(vccd2),
		.VSSD1(vssd2),

		.VSSD_PAD(vssd2_pad)

    	);

	// Instantiate analog pads in user area 1 using the custom analog pad
    	sky130_ef_io__analog_pad user1_analog_pad [ANALOG_PADS_1-2:0]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.P_PAD(mprj_io[19-2:19-ANALOG_PADS_1]),

		.P_CORE(mprj_analog[ANALOG_PADS_1-2:0])
    	);

	// Last analog pad is a power pad, to provide a clamp resource.
    	sky130_ef_io__top_power_hvc user1_analog_pad_with_clamp  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.P_PAD(mprj_io[19-1]),

		

	.DRN_HVC(mprj_clamp_high[0]),
	.SRC_BDY_HVC(mprj_clamp_low[0]),
		.P_CORE(mprj_analog[ANALOG_PADS_1-1])
    	);

	// Instantiate analog pads in user area 2 using the custom analog pad.
    	sky130_ef_io__analog_pad user2_analog_pad [ANALOG_PADS_2-3:0]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.P_PAD(mprj_io[19+ANALOG_PADS_2-1:19+2]),

		.P_CORE(mprj_analog[ANALOG_PADS_2+ANALOG_PADS_1-1:ANALOG_PADS_1+2])
    	);

	// Last two analog pads are power pads, to provide clamp resources.
    	sky130_ef_io__top_power_hvc user2_analog_pad_with_clamp [1:0] (

		.P_PAD(mprj_io[19+1:19]),

		
	.DRN_HVC(mprj_clamp_high[2:1]),
	.SRC_BDY_HVC(mprj_clamp_low[2:1]),
		.P_CORE(mprj_analog[5+1:ANALOG_PADS_1])
    	);

	wire [2:0] dm_all =
    		{gpio_mode1_core, gpio_mode1_core, gpio_mode0_core};
	wire[2:0] flash_io0_mode =
		{flash_io0_ieb_core, flash_io0_ieb_core, flash_io0_oeb_core};
	wire[2:0] flash_io1_mode =
		{flash_io1_ieb_core, flash_io1_ieb_core, flash_io1_oeb_core};

	wire [6:0] vccd_const_one;  // Constant value for management pins
	wire [6:0] vssd_const_zero; // Constant value for management pins

	constant_block constant_value_inst [6:0] (
            .vccd(vccd),
            .vssd(vssd),
            .one(vccd_const_one),
            .zero(vssd_const_zero)
	);

	// Management clock input pad
	
	wire loop_zero_clock;
	wire loop_one_clock;
	sky130_ef_io__gpiov2_pad_wrapped clock_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(clock),
	
		.OUT(vssd_const_zero[0]),
		.OE_N(vccd_const_one[0]),
		.HLD_H_N(loop_one_clock),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_clock),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_clock),
		.ENABLE_VDDIO(vccd_const_one[0]),
		.INP_DIS(por),
		.IB_MODE_SEL(vssd_const_zero[0]),
		.VTRIP_SEL(vssd_const_zero[0]),
		.SLOW(vssd_const_zero[0]),
		.HLD_OVR(vssd_const_zero[0]),
		.ANALOG_EN(vssd_const_zero[0]),
		.ANALOG_SEL(vssd_const_zero[0]),
		.ANALOG_POL(vssd_const_zero[0]),
		.DM({vssd_const_zero[0], vssd_const_zero[0], vccd_const_one[0]}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(clock_core),
		.IN_H(),
		.TIE_HI_ESD(loop_one_clock),
		.TIE_LO_ESD(loop_zero_clock) );

    	// Management GPIO pad
	
	wire loop_zero_gpio;
	wire loop_one_gpio;
	sky130_ef_io__gpiov2_pad_wrapped gpio_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(gpio),
	
		.OUT(gpio_out_core),
		.OE_N(gpio_outenb_core),
		.HLD_H_N(loop_one_gpio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_gpio),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_gpio),
		.ENABLE_VDDIO(vccd_const_one[1]),
		.INP_DIS(gpio_inenb_core),
		.IB_MODE_SEL(vssd_const_zero[1]),
		.VTRIP_SEL(vssd_const_zero[1]),
		.SLOW(vssd_const_zero[1]),
		.HLD_OVR(vssd_const_zero[1]),
		.ANALOG_EN(vssd_const_zero[1]),
		.ANALOG_SEL(vssd_const_zero[1]),
		.ANALOG_POL(vssd_const_zero[1]),
		.DM(dm_all),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(gpio_in_core),
		.IN_H(),
		.TIE_HI_ESD(loop_one_gpio),
		.TIE_LO_ESD(loop_zero_gpio) );

	// Management Flash SPI pads
	
	wire loop_zero_flash_io0;
	wire loop_one_flash_io0;
	sky130_ef_io__gpiov2_pad_wrapped flash_io0_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(flash_io0),
	
		.OUT(flash_io0_do_core),
		.OE_N(flash_io0_oeb_core),
		.HLD_H_N(loop_one_flash_io0),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_flash_io0),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_flash_io0),
		.ENABLE_VDDIO(vccd_const_one[2]),
		.INP_DIS(flash_io0_ieb_core),
		.IB_MODE_SEL(vssd_const_zero[2]),
		.VTRIP_SEL(vssd_const_zero[2]),
		.SLOW(vssd_const_zero[2]),
		.HLD_OVR(vssd_const_zero[2]),
		.ANALOG_EN(vssd_const_zero[2]),
		.ANALOG_SEL(vssd_const_zero[2]),
		.ANALOG_POL(vssd_const_zero[2]),
		.DM(flash_io0_mode),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(flash_io0_di_core),
		.IN_H(),
		.TIE_HI_ESD(loop_one_flash_io0),
		.TIE_LO_ESD(loop_zero_flash_io0) );
	
	wire loop_zero_flash_io1;
	wire loop_one_flash_io1;
	sky130_ef_io__gpiov2_pad_wrapped flash_io1_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(flash_io1),
	
		.OUT(flash_io1_do_core),
		.OE_N(flash_io1_oeb_core),
		.HLD_H_N(loop_one_flash_io1),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_flash_io1),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_flash_io1),
		.ENABLE_VDDIO(vccd_const_one[3]),
		.INP_DIS(flash_io1_ieb_core),
		.IB_MODE_SEL(vssd_const_zero[3]),
		.VTRIP_SEL(vssd_const_zero[3]),
		.SLOW(vssd_const_zero[3]),
		.HLD_OVR(vssd_const_zero[3]),
		.ANALOG_EN(vssd_const_zero[3]),
		.ANALOG_SEL(vssd_const_zero[3]),
		.ANALOG_POL(vssd_const_zero[3]),
		.DM(flash_io1_mode),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(flash_io1_di_core),
		.IN_H(),
		.TIE_HI_ESD(loop_one_flash_io1),
		.TIE_LO_ESD(loop_zero_flash_io1) );

	
	wire loop_zero_flash_csb;
	wire loop_one_flash_csb;
	sky130_ef_io__gpiov2_pad_wrapped flash_csb_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(flash_csb),
	
		.OUT(flash_csb_core),
		.OE_N(flash_csb_oeb_core),
		.HLD_H_N(loop_one_flash_csb),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_flash_csb),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_flash_csb),
		.ENABLE_VDDIO(vccd_const_one[4]),
		.INP_DIS(vssd_const_zero[4]),
		.IB_MODE_SEL(vssd_const_zero[4]),
		.VTRIP_SEL(vssd_const_zero[4]),
		.SLOW(vssd_const_zero[4]),
		.HLD_OVR(vssd_const_zero[4]),
		.ANALOG_EN(vssd_const_zero[4]),
		.ANALOG_SEL(vssd_const_zero[4]),
		.ANALOG_POL(vssd_const_zero[4]),
		.DM({vccd_const_one[4], vccd_const_one[4], vssd_const_zero[4]}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(),
		.IN_H(),
		.TIE_HI_ESD(loop_one_flash_csb),
		.TIE_LO_ESD(loop_zero_flash_csb));
	
	wire loop_zero_flash_clk;
	wire loop_one_flash_clk;
	sky130_ef_io__gpiov2_pad_wrapped flash_clk_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(flash_clk),
	
		.OUT(flash_clk_core),
		.OE_N(flash_clk_oeb_core),
		.HLD_H_N(loop_one_flash_clk),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_flash_clk),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_flash_clk),
		.ENABLE_VDDIO(vccd_const_one[5]),
		.INP_DIS(vssd_const_zero[5]),
		.IB_MODE_SEL(vssd_const_zero[5]),
		.VTRIP_SEL(vssd_const_zero[5]),
		.SLOW(vssd_const_zero[5]),
		.HLD_OVR(vssd_const_zero[5]),
		.ANALOG_EN(vssd_const_zero[5]),
		.ANALOG_SEL(vssd_const_zero[5]),
		.ANALOG_POL(vssd_const_zero[5]),
		.DM({vccd_const_one[5], vccd_const_one[5], vssd_const_zero[5]}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(),
		.IN_H(),
		.TIE_HI_ESD(loop_one_flash_clk),
		.TIE_LO_ESD(loop_zero_flash_clk));

	// NOTE:  The analog_out pad from the raven chip has been replaced by
    	// the digital reset input resetb on caravel due to the lack of an on-board
    	// power-on-reset circuit.  The XRES pad is used for providing a glitch-
    	// free reset.

	wire xresloop;
	wire xres_zero_loop;
	sky130_fd_io__top_xres4v2 resetb_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		
		    .PAD(resetb),
		
		.TIE_WEAK_HI_H(xresloop),   // Loop-back connection to pad through pad_a_esd_h
		.TIE_HI_ESD(),
		.TIE_LO_ESD(xres_zero_loop),
		.PAD_A_ESD_H(xresloop),
		.XRES_H_N(resetb_core_h),
		.DISABLE_PULLUP_H(xres_zero_loop),  // 0 = enable pull-up on reset pad
		.ENABLE_H(porb_h),	    	    // Power-on-reset
		.EN_VDDIO_SIG_H(xres_zero_loop),    // No idea.
		.INP_SEL_H(xres_zero_loop),	    // 1 = use filt_in_h else filter the pad input
		.FILT_IN_H(xres_zero_loop),	    // Alternate input for glitch filter
		.PULLUP_H(xres_zero_loop),	    // Pullup connection for alternate filter input
		.ENABLE_VDDIO(vccd_const_one[6])
    	);

	// Corner cells (These are overlay cells;  it is not clear what is normally
    	// supposed to go under them.)

	    sky130_ef_io__corner_pad mgmt_corner [1:0] (

		.VSSIO(vssio),
		.VDDIO(vddio),
		.VDDIO_Q(vddio_q),
		.VSSIO_Q(vssio_q),
		.AMUXBUS_A(analog_a),
		.AMUXBUS_B(analog_b),
		.VSSD(vssd),
		.VSSA(vssa),
		.VSWITCH(vddio),
		.VDDA(vdda),
		.VCCD(vccd),
		.VCCHIB(vccd)

    	    );

	    sky130_ef_io__corner_pad user1_corner (

		.VSSIO(vssio),
		.VDDIO(vddio),
		.VDDIO_Q(vddio_q),
		.VSSIO_Q(vssio_q),
		.AMUXBUS_A(analog_a),
		.AMUXBUS_B(analog_b),
		.VSSD(vssd),
		.VSSA(vssa1),
		.VSWITCH(vddio),
		.VDDA(vdda1),
		.VCCD(vccd),
		.VCCHIB(vccd)

    	    );
	    sky130_ef_io__corner_pad user2_corner (

		.VSSIO(vssio),
		.VDDIO(vddio),
		.VDDIO_Q(vddio_q),
		.VSSIO_Q(vssio_q),
		.AMUXBUS_A(analog_a),
		.AMUXBUS_B(analog_b),
		.VSSD(vssd),
		.VSSA(vssa2),
		.VSWITCH(vddio),
		.VDDA(vdda2),
		.VCCD(vccd),
		.VCCHIB(vccd)

    	    );

	mprj_io #(
		.AREA1PADS(19 - ANALOG_PADS_1),
		.TOTAL_PADS((19 + 19) - ANALOG_PADS_1 - ANALOG_PADS_2)
	) mprj_pads (
		.vddio(vddio),
		.vssio(vssio),
		.vccd(vccd),
		.vssd(vssd),
		.vdda1(vdda1),
		.vdda2(vdda2),
		.vssa1(vssa1),
		.vssa2(vssa2),
		.vddio_q(vddio_q),
		.vssio_q(vssio_q),
		.analog_a(analog_a),
		.analog_b(analog_b),
		.porb_h(porb_h),
		.vccd_conb(mprj_io_one),

		.io({mprj_io[(19 + 19)-1:19+ANALOG_PADS_2],
			     mprj_io[19-ANALOG_PADS_1-1:0]}),
		.io_out(mprj_io_out),
		.oeb(mprj_io_oeb),
		.enh(mprj_io_enh),
		.inp_dis(mprj_io_inp_dis),
		.ib_mode_sel(mprj_io_ib_mode_sel),
		.vtrip_sel(mprj_io_vtrip_sel),
		.holdover(mprj_io_holdover),
		.slow_sel(mprj_io_slow_sel),
		.analog_en(mprj_io_analog_en),
		.analog_sel(mprj_io_analog_sel),
		.analog_pol(mprj_io_analog_pol),
		.dm(mprj_io_dm),
		.io_in(mprj_io_in),
		.io_in_3v3(mprj_io_in_3v3),
		.analog_io(mprj_gpio_analog),
		.analog_noesd_io(mprj_gpio_noesd)
	);

endmodule
// `default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// `default_nettype none
module chip_io(
	// Package Pins
	inout  vddio_pad,		// Common padframe/ESD supply
	inout  vddio_pad2,
	inout  vssio_pad,		// Common padframe/ESD ground
	inout  vssio_pad2,
	inout  vccd_pad,		// Common 1.8V supply
	inout  vssd_pad,		// Common digital ground
	inout  vdda_pad,		// Management analog 3.3V supply
	inout  vssa_pad,		// Management analog ground
	inout  vdda1_pad,		// User area 1 3.3V supply
	inout  vdda1_pad2,		
	inout  vdda2_pad,		// User area 2 3.3V supply
	inout  vssa1_pad,		// User area 1 analog ground
	inout  vssa1_pad2,
	inout  vssa2_pad,		// User area 2 analog ground
	inout  vccd1_pad,		// User area 1 1.8V supply
	inout  vccd2_pad,		// User area 2 1.8V supply
	inout  vssd1_pad,		// User area 1 digital ground
	inout  vssd2_pad,		// User area 2 digital ground

	// Core Side
	inout  vddio,		// Common padframe/ESD supply
	inout  vssio,		// Common padframe/ESD ground
	inout  vccd,		// Common 1.8V supply
	inout  vssd,		// Common digital ground
	inout  vdda,		// Management analog 3.3V supply
	inout  vssa,		// Management analog ground
	inout  vdda1,		// User area 1 3.3V supply
	inout  vdda2,		// User area 2 3.3V supply
	inout  vssa1,		// User area 1 analog ground
	inout  vssa2,		// User area 2 analog ground
	inout  vccd1,		// User area 1 1.8V supply
	inout  vccd2,		// User area 2 1.8V supply
	inout  vssd1,		// User area 1 digital ground
	inout  vssd2,		// User area 2 digital ground

	inout  gpio,
	input  clock,
	input  resetb,
	output flash_csb,
	output flash_clk,
	inout  flash_io0,
	inout  flash_io1,
	// Chip Core Interface
	input  porb_h,
	input  por,
	output resetb_core_h,
	output clock_core,
	input  gpio_out_core,
	output gpio_in_core,
	input  gpio_mode0_core,
	input  gpio_mode1_core,
	input  gpio_outenb_core,
	input  gpio_inenb_core,
	input  flash_csb_core,
	input  flash_clk_core,
	input  flash_csb_oeb_core,
	input  flash_clk_oeb_core,
	input  flash_io0_oeb_core,
	input  flash_io1_oeb_core,
	input  flash_io0_ieb_core,
	input  flash_io1_ieb_core,
	input  flash_io0_do_core,
	input  flash_io1_do_core,
	output flash_io0_di_core,
	output flash_io1_di_core,
	// User project IOs
	inout [(19 + 19)-1:0] mprj_io,
	input [(19 + 19)-1:0] mprj_io_out,
	input [(19 + 19)-1:0] mprj_io_oeb,
	input [(19 + 19)-1:0] mprj_io_inp_dis,
	input [(19 + 19)-1:0] mprj_io_ib_mode_sel,
	input [(19 + 19)-1:0] mprj_io_vtrip_sel,
	input [(19 + 19)-1:0] mprj_io_slow_sel,
	input [(19 + 19)-1:0] mprj_io_holdover,
	input [(19 + 19)-1:0] mprj_io_analog_en,
	input [(19 + 19)-1:0] mprj_io_analog_sel,
	input [(19 + 19)-1:0] mprj_io_analog_pol,
	input [(19 + 19)*3-1:0] mprj_io_dm,
	output [(19 + 19)-1:0] mprj_io_in,
	// Loopbacks to constant value 1 in the 1.8V domain
	input [(19 + 19)-1:0] mprj_io_one,
	// User project direct access to gpio pad connections for analog
	// (all but the lowest-numbered 7 pads)
	inout [(19 + 19)-10:0] mprj_analog_io
);

    // To be considered:  Master hold signal on all user pads (?)
    // For now, set holdh_n to 1 internally (NOTE:  This is in the
    // VDDIO 3.3V domain)
    // and setting enh to porb_h.

    wire [(19 + 19)-1:0] mprj_io_enh;

    assign mprj_io_enh = {(19 + 19){porb_h}};
	
	wire analog_a, analog_b;
	wire vddio_q, vssio_q;

	// Instantiate power and ground pads for management domain
	// 12 pads:  vddio, vssio, vdda, vssa, vccd, vssd
	// One each HV and LV clamp.

	// HV clamps connect between one HV power rail and one ground
	// LV clamps have two clamps connecting between any two LV power
	// rails and grounds, and one back-to-back diode which connects
	// between the first LV clamp ground and any other ground.

    	sky130_ef_io__vddio_hvc_clamped_pad \mgmt_vddio_hvclamp_pad[0]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDIO_PAD(vddio_pad)

    	);

	// lies in user area 2
    	sky130_ef_io__vddio_hvc_clamped_pad \mgmt_vddio_hvclamp_pad[1]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDIO_PAD(vddio_pad2)

    	);

    	sky130_ef_io__vdda_hvc_clamped_pad mgmt_vdda_hvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDA_PAD(vdda_pad)

    	);

    	sky130_ef_io__vccd_lvc_clamped_pad mgmt_vccd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VCCD_PAD(vccd_pad)

    	);

    	sky130_ef_io__vssio_hvc_clamped_pad \mgmt_vssio_hvclamp_pad[0]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSIO_PAD(vssio_pad)

    	);

    	sky130_ef_io__vssio_hvc_clamped_pad \mgmt_vssio_hvclamp_pad[1]  (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSIO_PAD(vssio_pad2)

    	);

    	sky130_ef_io__vssa_hvc_clamped_pad mgmt_vssa_hvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSA_PAD(vssa_pad)

    	);

    	sky130_ef_io__vssd_lvc_clamped_pad mgmt_vssd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSD_PAD(vssd_pad)

    	);

	// Instantiate power and ground pads for user 1 domain
	// 8 pads:  vdda, vssa, vccd, vssd;  One each HV and LV clamp.

    	sky130_ef_io__vdda_hvc_clamped_pad \user1_vdda_hvclamp_pad[0] (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDA_PAD(vdda1_pad)

    	);

		sky130_ef_io__vdda_hvc_clamped_pad \user1_vdda_hvclamp_pad[1] (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDA_PAD(vdda1_pad2)

    	);

    	sky130_ef_io__vccd_lvc_clamped3_pad user1_vccd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		.VCCD1(vccd1),
		.VSSD1(vssd1),

		.VCCD_PAD(vccd1_pad)

    	);

    	sky130_ef_io__vssa_hvc_clamped_pad \user1_vssa_hvclamp_pad[0] (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSA_PAD(vssa1_pad)

    	);


    	sky130_ef_io__vssa_hvc_clamped_pad \user1_vssa_hvclamp_pad[1] (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSA_PAD(vssa1_pad2)

    	);

    	sky130_ef_io__vssd_lvc_clamped3_pad user1_vssd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa1),
	.VDDA(vdda1),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		.VCCD1(vccd1),
		.VSSD1(vssd1),

		.VSSD_PAD(vssd1_pad)

    	);

	// Instantiate power and ground pads for user 2 domain
	// 8 pads:  vdda, vssa, vccd, vssd;  One each HV and LV clamp.

    	sky130_ef_io__vdda_hvc_clamped_pad user2_vdda_hvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VDDA_PAD(vdda2_pad)

    	);

    	sky130_ef_io__vccd_lvc_clamped3_pad user2_vccd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		.VCCD1(vccd2),
		.VSSD1(vssd2),

		.VCCD_PAD(vccd2_pad)

    	);

    	sky130_ef_io__vssa_hvc_clamped_pad user2_vssa_hvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),

		.VSSA_PAD(vssa2_pad)

    	);

    	sky130_ef_io__vssd_lvc_clamped3_pad user2_vssd_lvclamp_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa2),
	.VDDA(vdda2),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		.VCCD1(vccd2),
		.VSSD1(vssd2),

		.VSSD_PAD(vssd2_pad)

    	);

	wire [2:0] dm_all =
    		{gpio_mode1_core, gpio_mode1_core, gpio_mode0_core};
	wire[2:0] flash_io0_mode =
		{flash_io0_ieb_core, flash_io0_ieb_core, flash_io0_oeb_core};
	wire[2:0] flash_io1_mode =
		{flash_io1_ieb_core, flash_io1_ieb_core, flash_io1_oeb_core};

    wire [6:0] vccd_const_one;	// Constant value for management pins
    wire [6:0] vssd_const_zero;	// Constant value for management pins

    constant_block constant_value_inst [6:0] (
	.vccd(vccd),
	.vssd(vssd),
	.one(vccd_const_one),
	.zero(vssd_const_zero)
    );

	// Management clock input pad
	
	wire loop_zero_clock;
	wire loop_one_clock;
	sky130_ef_io__gpiov2_pad_wrapped clock_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(clock),
	
		.OUT(vssd_const_zero[0]),
		.OE_N(vccd_const_one[0]),
		.HLD_H_N(loop_one_clock),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_clock),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_clock),
		.ENABLE_VDDIO(vccd_const_one[0]),
		.INP_DIS(por),
		.IB_MODE_SEL(vssd_const_zero[0]),
		.VTRIP_SEL(vssd_const_zero[0]),
		.SLOW(vssd_const_zero[0]),
		.HLD_OVR(vssd_const_zero[0]),
		.ANALOG_EN(vssd_const_zero[0]),
		.ANALOG_SEL(vssd_const_zero[0]),
		.ANALOG_POL(vssd_const_zero[0]),
		.DM({vssd_const_zero[0], vssd_const_zero[0], vccd_const_one[0]}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(clock_core),
		.IN_H(),
		.TIE_HI_ESD(loop_one_clock),
		.TIE_LO_ESD(loop_zero_clock) );

    // Management GPIO pad
	
	wire loop_zero_gpio;
	wire loop_one_gpio;
	sky130_ef_io__gpiov2_pad_wrapped gpio_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(gpio),
	
		.OUT(gpio_out_core),
		.OE_N(gpio_outenb_core),
		.HLD_H_N(loop_one_gpio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_gpio),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_gpio),
		.ENABLE_VDDIO(vccd_const_one[1]),
		.INP_DIS(gpio_inenb_core),
		.IB_MODE_SEL(vssd_const_zero[1]),
		.VTRIP_SEL(vssd_const_zero[1]),
		.SLOW(vssd_const_zero[1]),
		.HLD_OVR(vssd_const_zero[1]),
		.ANALOG_EN(vssd_const_zero[1]),
		.ANALOG_SEL(vssd_const_zero[1]),
		.ANALOG_POL(vssd_const_zero[1]),
		.DM(dm_all),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(gpio_in_core),
		.IN_H(),
		.TIE_HI_ESD(loop_one_gpio),
		.TIE_LO_ESD(loop_zero_gpio) );

	// Management Flash SPI pads
	
	wire loop_zero_flash_io0;
	wire loop_one_flash_io0;
	sky130_ef_io__gpiov2_pad_wrapped flash_io0_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(flash_io0),
	
		.OUT(flash_io0_do_core),
		.OE_N(flash_io0_oeb_core),
		.HLD_H_N(loop_one_flash_io0),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_flash_io0),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_flash_io0),
		.ENABLE_VDDIO(vccd_const_one[2]),
		.INP_DIS(flash_io0_ieb_core),
		.IB_MODE_SEL(vssd_const_zero[2]),
		.VTRIP_SEL(vssd_const_zero[2]),
		.SLOW(vssd_const_zero[2]),
		.HLD_OVR(vssd_const_zero[2]),
		.ANALOG_EN(vssd_const_zero[2]),
		.ANALOG_SEL(vssd_const_zero[2]),
		.ANALOG_POL(vssd_const_zero[2]),
		.DM(flash_io0_mode),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(flash_io0_di_core),
		.IN_H(),
		.TIE_HI_ESD(loop_one_flash_io0),
		.TIE_LO_ESD(loop_zero_flash_io0) );
	
	
	wire loop_zero_flash_io1;
	wire loop_one_flash_io1;
	sky130_ef_io__gpiov2_pad_wrapped flash_io1_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(flash_io1),
	
		.OUT(flash_io1_do_core),
		.OE_N(flash_io1_oeb_core),
		.HLD_H_N(loop_one_flash_io1),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_flash_io1),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_flash_io1),
		.ENABLE_VDDIO(vccd_const_one[3]),
		.INP_DIS(flash_io1_ieb_core),
		.IB_MODE_SEL(vssd_const_zero[3]),
		.VTRIP_SEL(vssd_const_zero[3]),
		.SLOW(vssd_const_zero[3]),
		.HLD_OVR(vssd_const_zero[3]),
		.ANALOG_EN(vssd_const_zero[3]),
		.ANALOG_SEL(vssd_const_zero[3]),
		.ANALOG_POL(vssd_const_zero[3]),
		.DM(flash_io1_mode),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(flash_io1_di_core),
		.IN_H(),
		.TIE_HI_ESD(loop_one_flash_io1),
		.TIE_LO_ESD(loop_zero_flash_io1) );

	
	wire loop_zero_flash_csb;
	wire loop_one_flash_csb;
	sky130_ef_io__gpiov2_pad_wrapped flash_csb_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(flash_csb),
	
		.OUT(flash_csb_core),
		.OE_N(flash_csb_oeb_core),
		.HLD_H_N(loop_one_flash_csb),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_flash_csb),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_flash_csb),
		.ENABLE_VDDIO(vccd_const_one[4]),
		.INP_DIS(vssd_const_zero[4]),
		.IB_MODE_SEL(vssd_const_zero[4]),
		.VTRIP_SEL(vssd_const_zero[4]),
		.SLOW(vssd_const_zero[4]),
		.HLD_OVR(vssd_const_zero[4]),
		.ANALOG_EN(vssd_const_zero[4]),
		.ANALOG_SEL(vssd_const_zero[4]),
		.ANALOG_POL(vssd_const_zero[4]),
		.DM({vccd_const_one[4], vccd_const_one[4], vssd_const_zero[4]}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(),
		.IN_H(),
		.TIE_HI_ESD(loop_one_flash_csb),
		.TIE_LO_ESD(loop_zero_flash_csb));
	
	wire loop_zero_flash_clk;
	wire loop_one_flash_clk;
	sky130_ef_io__gpiov2_pad_wrapped flash_clk_pad (
	
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
	
		.PAD(flash_clk),
	
		.OUT(flash_clk_core),
		.OE_N(flash_clk_oeb_core),
		.HLD_H_N(loop_one_flash_clk),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(loop_zero_flash_clk),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(loop_zero_flash_clk),
		.ENABLE_VDDIO(vccd_const_one[5]),
		.INP_DIS(vssd_const_zero[5]),
		.IB_MODE_SEL(vssd_const_zero[5]),
		.VTRIP_SEL(vssd_const_zero[5]),
		.SLOW(vssd_const_zero[5]),
		.HLD_OVR(vssd_const_zero[5]),
		.ANALOG_EN(vssd_const_zero[5]),
		.ANALOG_SEL(vssd_const_zero[5]),
		.ANALOG_POL(vssd_const_zero[5]),
		.DM({vccd_const_one[5], vccd_const_one[5], vssd_const_zero[5]}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(),
		.IN_H(),
		.TIE_HI_ESD(loop_one_flash_clk),
		.TIE_LO_ESD(loop_zero_flash_clk));

	// NOTE:  The analog_out pad from the raven chip has been replaced by
    	// the digital reset input resetb on caravel due to the lack of an on-board
    	// power-on-reset circuit.  The XRES pad is used for providing a glitch-
    	// free reset.

	wire xresloop;
	wire xres_vss_loop;
	sky130_fd_io__top_xres4v2 resetb_pad (
		
	.AMUXBUS_A(analog_a),
	.AMUXBUS_B(analog_b),
	.VSSA(vssa),
	.VDDA(vdda),
	.VSWITCH(vddio),
	.VDDIO_Q(vddio_q),
	.VCCHIB(vccd),
	.VDDIO(vddio),
	.VCCD(vccd),
	.VSSIO(vssio),
	.VSSD(vssd),
	.VSSIO_Q(vssio_q),
		
		    .PAD(resetb),
		
		.TIE_WEAK_HI_H(xresloop),   // Loop-back connection to pad through pad_a_esd_h
		.TIE_HI_ESD(),
		.TIE_LO_ESD(xres_vss_loop),
		.PAD_A_ESD_H(xresloop),
		.XRES_H_N(resetb_core_h),
		.DISABLE_PULLUP_H(xres_vss_loop), // 0 = enable pull-up on reset pad
		.ENABLE_H(porb_h),	 	  // Power-on-reset
   		.EN_VDDIO_SIG_H(xres_vss_loop),	  // No idea.
   		.INP_SEL_H(xres_vss_loop),	  // 1 = use filt_in_h else filter the pad input
   		.FILT_IN_H(xres_vss_loop),	  // Alternate input for glitch filter
   		.PULLUP_H(xres_vss_loop),	  // Pullup connection for alternate filter input
		.ENABLE_VDDIO(vccd_const_one[6])
    	);

	// Corner cells (These are overlay cells;  it is not clear what is normally
    	// supposed to go under them.)

	    sky130_ef_io__corner_pad mgmt_corner [1:0] (

		.VSSIO(vssio),
		.VDDIO(vddio),
		.VDDIO_Q(vddio_q),
		.VSSIO_Q(vssio_q),
		.AMUXBUS_A(analog_a),
		.AMUXBUS_B(analog_b),
		.VSSD(vssd),
		.VSSA(vssa),
		.VSWITCH(vddio),
		.VDDA(vdda),
		.VCCD(vccd),
		.VCCHIB(vccd)

    	    );
	    sky130_ef_io__corner_pad user1_corner (

		.VSSIO(vssio),
		.VDDIO(vddio),
		.VDDIO_Q(vddio_q),
		.VSSIO_Q(vssio_q),
		.AMUXBUS_A(analog_a),
		.AMUXBUS_B(analog_b),
		.VSSD(vssd),
		.VSSA(vssa1),
		.VSWITCH(vddio),
		.VDDA(vdda1),
		.VCCD(vccd),
		.VCCHIB(vccd)

    	    );
	    sky130_ef_io__corner_pad user2_corner (

		.VSSIO(vssio),
		.VDDIO(vddio),
		.VDDIO_Q(vddio_q),
		.VSSIO_Q(vssio_q),
		.AMUXBUS_A(analog_a),
		.AMUXBUS_B(analog_b),
		.VSSD(vssd),
		.VSSA(vssa2),
		.VSWITCH(vddio),
		.VDDA(vdda2),
		.VCCD(vccd),
		.VCCHIB(vccd)

    	    );

	mprj_io mprj_pads(
		.vddio(vddio),
		.vssio(vssio),
		.vccd(vccd),
		.vssd(vssd),
		.vdda1(vdda1),
		.vdda2(vdda2),
		.vssa1(vssa1),
		.vssa2(vssa2),
		.vddio_q(vddio_q),
		.vssio_q(vssio_q),
		.analog_a(analog_a),
		.analog_b(analog_b),
		.porb_h(porb_h),
		.vccd_conb(mprj_io_one),
		.io(mprj_io),
		.io_out(mprj_io_out),
		.oeb(mprj_io_oeb),
		.enh(mprj_io_enh),
		.inp_dis(mprj_io_inp_dis),
		.ib_mode_sel(mprj_io_ib_mode_sel),
		.vtrip_sel(mprj_io_vtrip_sel),
		.holdover(mprj_io_holdover),
		.slow_sel(mprj_io_slow_sel),
		.analog_en(mprj_io_analog_en),
		.analog_sel(mprj_io_analog_sel),
		.analog_pol(mprj_io_analog_pol),
		.dm(mprj_io_dm),
		.io_in(mprj_io_in),
		.analog_io(mprj_analog_io)
	);

endmodule
// `default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module mprj_logic_high (

    inout	   vccd1,
    inout	   vssd1,

    output [462:0] HI
);
sky130_fd_sc_hd__conb_1 insts [462:0] (

                .VPWR(vccd1),
                .VGND(vssd1),
                .VPB(vccd1),
                .VNB(vssd1),

                .HI(HI),
                .LO()
        );
endmodule
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module mprj2_logic_high (

    inout	   vccd2,
    inout	   vssd2,

    output         HI
);
sky130_fd_sc_hd__conb_1 inst (

                .VPWR(vccd2),
                .VGND(vssd2),
                .VPB(vccd2),
                .VNB(vssd2),

                .HI(HI),
                .LO()
        );
endmodule
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*----------------------------------------------------------------------*/
/* Buffers protecting the management region from the user region.	*/
/* This mainly consists of tristate buffers that are enabled by a	*/
/* "logic 1" output connected to the user's VCCD domain.  This ensures	*/
/* that the buffer is disabled and the output high-impedence when the	*/
/* user 1.8V supply is absent.						*/
/*----------------------------------------------------------------------*/
/* Because there is no tristate buffer with a non-inverted enable, a	*/
/* tristate inverter with non-inverted enable is used in series with	*/
/* another (normal) inverter.						*/
/*----------------------------------------------------------------------*/
/* For the sake of placement/routing, one conb (logic 1) cell is used	*/
/* for every buffer.							*/
/*----------------------------------------------------------------------*/
/* 10/3/2022:  Removed tri-state buffers in favor of AND gates;  i.e.,	*/
/* if the user project is powered down, then the outputs are grounded	*/
/* rather than tristated.  Other explicitly-referenced gates removed	*/
/* with the assumption that all outputs will be buffered as needed by	*/
/* the synthesis tools.  Therefore the only restrictions needed on the	*/
/* synthesis tools is the list of input signals that must not be	*/
/* buffered because they are allowed to be floating.			*/
/*----------------------------------------------------------------------*/

module mgmt_protect (

    inout	  vccd,
    inout	  vssd,
    inout	  vccd1,
    inout	  vssd1,
    inout	  vccd2,
    inout	  vssd2,
    inout	  vdda1,
    inout	  vssa1,
    inout	  vdda2,
    inout	  vssa2,


    input 	  caravel_clk,
    input 	  caravel_clk2,
    input	  caravel_rstn,
    input 	  mprj_cyc_o_core,
    input 	  mprj_stb_o_core,
    input         mprj_we_o_core,
    input [3:0]   mprj_sel_o_core,
    input [31:0]  mprj_adr_o_core,
    input [31:0]  mprj_dat_o_core,
    input [2:0]	  user_irq_core,

    output [31:0] mprj_dat_i_core,
    output	  mprj_ack_i_core,

    input  	  mprj_iena_wb,		// Enable wishbone from user project

    // All signal in/out directions are the reverse of the signal
    // names at the buffer intrface.

    output [127:0] la_data_in_mprj,
    input  [127:0] la_data_out_mprj,
    input  [127:0] la_oenb_mprj,
    input  [127:0] la_iena_mprj,

    input  [127:0] la_data_out_core,
    output [127:0] la_data_in_core,
    output [127:0] la_oenb_core,

    input  [2:0]  user_irq_ena,

    output 	  user_clock,
    output 	  user_clock2,
    output 	  user_reset,
    output 	  mprj_cyc_o_user,
    output 	  mprj_stb_o_user,
    output 	  mprj_we_o_user,
    output [3:0]  mprj_sel_o_user,
    output [31:0] mprj_adr_o_user,
    output [31:0] mprj_dat_o_user,
    input  [31:0] mprj_dat_i_user,
    input	  mprj_ack_i_user,
    output [2:0]  user_irq,
    output	  user1_vcc_powergood,
    output	  user2_vcc_powergood,
    output	  user1_vdd_powergood,
    output	  user2_vdd_powergood
);

	wire [462:0] mprj_logic1;
	wire	     mprj2_logic1;

	wire mprj_vdd_logic1_h;
	wire mprj2_vdd_logic1_h;
	wire mprj_vdd_logic1;
	wire mprj2_vdd_logic1;


	wire [127:0] la_data_in_mprj_bar;
	wire [2:0] user_irq_bar;

	wire [127:0] la_data_in_enable;
	wire [127:0] la_data_out_enable;
	wire [2:0] user_irq_enable;
	wire 	   wb_in_enable;

	wire [31:0] mprj_dat_i_core_bar;
	wire 	    mprj_ack_i_core_bar;

        mprj_logic_high mprj_logic_high_inst (

                .vccd1(vccd1),
                .vssd1(vssd1),

                .HI(mprj_logic1)
        );

        mprj2_logic_high mprj2_logic_high_inst (

                .vccd2(vccd2),
                .vssd2(vssd2),

                .HI(mprj2_logic1)
        );

	// Logic high in the VDDA (3.3V) domains

	mgmt_protect_hv powergood_check (

	    .vccd(vccd),
	    .vssd(vssd),
	    .vdda1(vdda1),
	    .vssa1(vssa1),
	    .vdda2(vdda2),
	    .vssa2(vssa2),

	    .mprj_vdd_logic1(mprj_vdd_logic1),
	    .mprj2_vdd_logic1(mprj2_vdd_logic1)
	);

	// Buffering from the user side to the management side.
	// NOTE:  This is intended to be better protected, by a full
	// chain of an lv-to-hv buffer followed by an hv-to-lv buffer.
	// This serves as a placeholder until that configuration is
	// checked and characterized.  The function below forces the
	// data input to the management core to be a solid logic 0 when
	// the user project is powered down.

	assign la_data_in_enable = la_iena_mprj & mprj_logic1[457:330];

	sky130_fd_sc_hd__nand2_4 user_to_mprj_in_gates [127:0] (

                .VPWR(vccd),
                .VGND(vssd),
                .VPB(vccd),
                .VNB(vssd),

		.Y(la_data_in_mprj_bar),
		.A(la_data_out_core),		// may be floating
		.B(la_data_in_enable)
	);

	assign la_data_in_mprj = ~la_data_in_mprj_bar;

	// Protection, similar to the above, for the three user IRQ lines

	assign user_irq_enable = user_irq_ena & mprj_logic1[460:458];

	sky130_fd_sc_hd__nand2_4 user_irq_gates [2:0] (

                .VPWR(vccd),
                .VGND(vssd),
                .VPB(vccd),
                .VNB(vssd),

		.Y(user_irq_bar),
		.A(user_irq_core),		// may be floating
		.B(user_irq_enable)
	);

	assign user_irq = ~user_irq_bar;

	// Protection, similar to the above, for the return
	// signals from user area to managment on the wishbone bus

	assign wb_in_enable = mprj_iena_wb & mprj_logic1[462];

	sky130_fd_sc_hd__nand2_4 user_wb_dat_gates [31:0] (

                .VPWR(vccd),
                .VGND(vssd),
                .VPB(vccd),
                .VNB(vssd),

		.Y(mprj_dat_i_core_bar),
		.A(mprj_dat_i_user),		// may be floating
		.B(wb_in_enable)
	);

	assign mprj_dat_i_core = ~mprj_dat_i_core_bar;

	sky130_fd_sc_hd__nand2_4 user_wb_ack_gate (

                .VPWR(vccd),
                .VGND(vssd),
                .VPB(vccd),
                .VNB(vssd),

		.Y(mprj_ack_i_core_bar),
		.A(mprj_ack_i_user),		// may be floating
		.B(wb_in_enable)
	);

	assign mprj_ack_i_core = ~mprj_ack_i_core_bar;

	// The remaining circuitry guards against the management
	// SoC dumping current into the user project area when
	// the user project area is powered down.
	
	assign user_reset      = (~caravel_rstn) & mprj_logic1[0];
	assign user_clock      = caravel_clk     & mprj_logic1[1];
	assign user_clock2     = caravel_clk2    & mprj_logic1[2];
	assign mprj_cyc_o_user = mprj_cyc_o_core & mprj_logic1[3];
	assign mprj_stb_o_user = mprj_stb_o_core & mprj_logic1[4];
	assign mprj_we_o_user  = mprj_we_o_core  & mprj_logic1[5];
	assign mprj_sel_o_user = mprj_sel_o_core & mprj_logic1[9:6];
	assign mprj_adr_o_user = mprj_adr_o_core & mprj_logic1[41:10];
	assign mprj_dat_o_user = mprj_dat_o_core & mprj_logic1[73:42];

	/* Project data out from the managment side to the user project	*/
	/* area when the user project is powered down.			*/

	assign la_data_out_enable = (~la_oenb_mprj) & mprj_logic1[201:74];
	assign la_data_in_core = la_data_out_mprj & la_data_out_enable;

	/* Project data out enable (bar) from the managment side to the	*/
	/* user project	area when the user project is powered down.	*/

	assign la_oenb_core = la_oenb_mprj & mprj_logic1[329:202];

	/* The conb cell output is a resistive connection directly to	*/
	/* the power supply, so when returning the user1_powergood	*/
	/* signal, make sure that it is buffered properly.		*/

	assign user1_vcc_powergood = mprj_logic1[461];
	assign user2_vcc_powergood = mprj2_logic1;
	assign user1_vdd_powergood = mprj_vdd_logic1;
	assign user2_vdd_powergood = mprj2_vdd_logic1;

endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*----------------------------------------------------------------------*/
/* mgmt_protect_hv:							*/
/*									*/
/* High voltage (3.3V) part of the mgmt_protect module.  Split out into	*/
/* a separate module and file so that the synthesis tools can handle it	*/
/* separately from the rest, since it uses a different standard cell	*/
/* library.  See the file mgmt_protect.v for a full description of the	*/
/* whole management protection method.					*/
/*----------------------------------------------------------------------*/

module mgmt_protect_hv (

    inout	vccd,
    inout	vssd,
    inout	vdda1,
    inout	vssa1,
    inout	vdda2,
    inout	vssa2,


    output	mprj_vdd_logic1,
    output	mprj2_vdd_logic1

);

    wire mprj_vdd_logic1_h;
    wire mprj2_vdd_logic1_h;


    // This is to emulate the substrate shorting grounds together for LVS
    // purposes
    assign vssa2 = vssa1;
    assign vssa1 = vssd;


    // Logic high in the VDDA (3.3V) domains

    sky130_fd_sc_hvl__conb_1 mprj_logic_high_hvl (

        .VPWR(vdda1),
        .VGND(vssa1),
        .VPB(vdda1),
        .VNB(vssa1),

        .HI(mprj_vdd_logic1_h),
        .LO()
    );

    sky130_fd_sc_hvl__conb_1 mprj2_logic_high_hvl (

        .VPWR(vdda2),
        .VGND(vssa2),
        .VPB(vdda2),
        .VNB(vssa2),

        .HI(mprj2_vdd_logic1_h),
        .LO()
    );

    // Level shift the logic high signals into the 1.8V domain

    sky130_fd_sc_hvl__lsbufhv2lv_1 mprj_logic_high_lv (

	.VPWR(vdda1),
	.VGND(vssd),
	.LVPWR(vccd),
	.VPB(vdda1),
	.VNB(vssd),

	.X(mprj_vdd_logic1),
	.A(mprj_vdd_logic1_h)
    );

    sky130_fd_sc_hvl__lsbufhv2lv_1 mprj2_logic_high_lv (

	.VPWR(vdda2),
	.VGND(vssd),
	.LVPWR(vccd),
	.VPB(vdda2),
	.VNB(vssd),

	.X(mprj2_vdd_logic1),
	.A(mprj2_vdd_logic1_h)
    );
endmodule

`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/* 
 *---------------------------------------------------------------------
 * See gpio_control_block for description.  This module is like
 * gpio_contro_block except that it has an additional two management-
 * Soc-facing pins, which are the out_enb line and the output line.
 * If the chip is configured for output with the oeb control
 * register = 1, then the oeb line is controlled by the additional
 * signal from the management SoC.  If the oeb control register = 0,
 * then the output is disabled completely.  The "io" line is input
 * only in this module.
 *
 *---------------------------------------------------------------------
 */

/*
 *---------------------------------------------------------------------
 *
 * This module instantiates a shift register chain that passes through
 * each gpio cell.  These are connected end-to-end around the padframe
 * periphery.  The purpose is to avoid a massive number of control
 * wires between the digital core and I/O, passing through the user area.
 *
 * See mprj_ctrl.v for the module that registers the data for each
 * I/O and drives the input to the shift register.
 *
 * Modified 7/24/2022 by Tim Edwards
 * Replaced the data delay with a negative edge-triggered flop
 * so that the serial data bit out from the module only changes on
 * the clock half cycle.  This avoids the need to fine-tune the clock
 * skew between GPIO blocks.
 *
 * Modified 10/05/2022 by Tim Edwards
 *
 *---------------------------------------------------------------------
 */

module gpio_control_block #(
    parameter PAD_CTRL_BITS = 13
) (
    
         inout vccd,
         inout vssd,
         inout vccd1,
         inout vssd1,
    

    // Power-on defaults
    input [PAD_CTRL_BITS-1:0] gpio_defaults,

    // Management Soc-facing signals
    input  	 resetn,		// Global reset, locally propagated
    output       resetn_out,
    input  	 serial_clock,		// Global clock, locally propatated
    output  	 serial_clock_out,
    input	 serial_load,		// Register load strobe
    output	 serial_load_out,

    output       mgmt_gpio_in,		// Management from pad (input only)
    input        mgmt_gpio_out,		// Management to pad (output only)
    input        mgmt_gpio_oeb,		// Management to pad (output only)

    // Serial data chain for pad configuration
    input  	 serial_data_in,
    output reg   serial_data_out,

    // User-facing signals
    input        user_gpio_out,		// User space to pad
    input        user_gpio_oeb,		// Output enable (user)
    output	 user_gpio_in,		// Pad to user space

    // Pad-facing signals (Pad GPIOv2)
    output	 pad_gpio_holdover,
    output	 pad_gpio_slow_sel,
    output	 pad_gpio_vtrip_sel,
    output       pad_gpio_inenb,
    output       pad_gpio_ib_mode_sel,
    output	 pad_gpio_ana_en,
    output	 pad_gpio_ana_sel,
    output	 pad_gpio_ana_pol,
    output [2:0] pad_gpio_dm,
    output       pad_gpio_outenb,
    output	 pad_gpio_out,
    input	 pad_gpio_in,

    // to provide a way to automatically disable/enable output
    // from the outside with needing a conb cell
    output	 one,
    output	 zero
);

    /* Parameters defining the bit offset of each function in the chain */
    localparam MGMT_EN = 0;
    localparam OEB = 1;
    localparam HLDH = 2;
    localparam INP_DIS = 3;
    localparam MOD_SEL = 4;
    localparam AN_EN = 5;
    localparam AN_SEL = 6;
    localparam AN_POL = 7;
    localparam SLOW = 8;
    localparam TRIP = 9;
    localparam DM = 10;

    /* Internally registered signals */
    reg	 	mgmt_ena;		// Enable management SoC to access pad
    reg	 	gpio_holdover;
    reg	 	gpio_slow_sel;
    reg	  	gpio_vtrip_sel;
    reg  	gpio_inenb;
    reg	 	gpio_ib_mode_sel;
    reg  	gpio_outenb;
    reg [2:0] 	gpio_dm;
    reg	 	gpio_ana_en;
    reg	 	gpio_ana_sel;
    reg	 	gpio_ana_pol;

    wire	one_unbuf;
    wire	zero_unbuf;

    wire gpio_logic1;

    /* Serial shift for the above (latched) values */
    reg [PAD_CTRL_BITS-1:0] shift_register;

    /* Latch the output on the clock negative edge */
    always @(negedge serial_clock or negedge resetn) begin
	if (resetn == 1'b0) begin
	    /* Clear the shift register output */
	    serial_data_out <= 1'b0;
        end else begin
	    serial_data_out <= shift_register[PAD_CTRL_BITS-1];
	end
    end

    /* Propagate the clock and reset signals so that they aren't wired	*/
    /* all over the chip, but are just wired between the blocks.	*/
    (* keep *) sky130_fd_sc_hd__clkbuf_8 BUF[2:0] (
    
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
    
        .A({serial_clock, resetn, serial_load}),
        .X({serial_clock_out, resetn_out, serial_load_out})
    );

    always @(posedge serial_clock or negedge resetn) begin
	if (resetn == 1'b0) begin
	    /* Clear shift register */
	    shift_register <= 'd0;
	end else begin
	    /* Shift data in */
	    shift_register <= {shift_register[PAD_CTRL_BITS-2:0], serial_data_in};
	end
    end

    always @(posedge serial_load or negedge resetn) begin
	if (resetn == 1'b0) begin
	    /* Initial state on reset depends on applied defaults */
	    mgmt_ena <= gpio_defaults[MGMT_EN];
	    gpio_holdover <= gpio_defaults[HLDH];
	    gpio_slow_sel <= gpio_defaults[SLOW];
	    gpio_vtrip_sel <= gpio_defaults[TRIP];
            gpio_ib_mode_sel <= gpio_defaults[MOD_SEL];
	    gpio_inenb <= gpio_defaults[INP_DIS];
	    gpio_outenb <= gpio_defaults[OEB];
	    gpio_dm <= gpio_defaults[DM+2:DM];
	    gpio_ana_en <= gpio_defaults[AN_EN];
	    gpio_ana_sel <= gpio_defaults[AN_SEL];
	    gpio_ana_pol <= gpio_defaults[AN_POL];
	end else begin
	    /* Load data */
	    mgmt_ena 	     <= shift_register[MGMT_EN];
	    gpio_outenb      <= shift_register[OEB];
	    gpio_holdover    <= shift_register[HLDH]; 
	    gpio_inenb 	     <= shift_register[INP_DIS];
	    gpio_ib_mode_sel <= shift_register[MOD_SEL];
	    gpio_ana_en      <= shift_register[AN_EN];
	    gpio_ana_sel     <= shift_register[AN_SEL];
	    gpio_ana_pol     <= shift_register[AN_POL];
	    gpio_slow_sel    <= shift_register[SLOW];
	    gpio_vtrip_sel   <= shift_register[TRIP];
	    gpio_dm 	     <= shift_register[DM+2:DM];

	end
    end

    /* These pad configuration signals are static and do not change	*/
    /* after setup.							*/

    assign pad_gpio_holdover 	= gpio_holdover;
    assign pad_gpio_slow_sel 	= gpio_slow_sel;
    assign pad_gpio_vtrip_sel	= gpio_vtrip_sel;
    assign pad_gpio_ib_mode_sel	= gpio_ib_mode_sel;
    assign pad_gpio_ana_en	= gpio_ana_en;
    assign pad_gpio_ana_sel	= gpio_ana_sel;
    assign pad_gpio_ana_pol	= gpio_ana_pol;
    assign pad_gpio_dm		= gpio_dm;
    assign pad_gpio_inenb 	= gpio_inenb;

    /* Implement pad control behavior depending on state of mgmt_ena */

    /* The pad value always goes back to the housekeeping module	*/

    assign mgmt_gpio_in = pad_gpio_in;

    /* For 2-wire interfaces, the mgmt_gpio_oeb line is tied high at	*/
    /* the control block.  In this case, the output enable state is	*/
    /* determined by the OEB configuration bit.				*/

    assign pad_gpio_outenb = (mgmt_ena) ? ((mgmt_gpio_oeb == 1'b1) ?
			gpio_outenb : 1'b0) : user_gpio_oeb;

    /* For 2-wire interfaces, if the pad is configured for pull-up or	*/
    /* pull-down, drive the output value locally to achieve the		*/
    /* expected pull.							*/

    assign pad_gpio_out = (mgmt_ena) ? ((mgmt_gpio_oeb == 1'b1) ?
			((gpio_dm[2:1] == 2'b01) ? ~gpio_dm[0] : mgmt_gpio_out) :
			mgmt_gpio_out) : user_gpio_out; 

    /* Buffer user_gpio_in with an enable that is set by the user domain vccd */

    gpio_logic_high gpio_logic_high (

            .vccd1(vccd1),
            .vssd1(vssd1),

            .gpio_logic1(gpio_logic1)
    );

    /* If user project area is powered down, zero the pad input value	*/
    /* going to the user project.					*/
    assign user_gpio_in = pad_gpio_in & gpio_logic1;

    (* keep *)
    sky130_fd_sc_hd__macro_sparecell spare_cell (

            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd)

    );

    sky130_fd_sc_hd__conb_1 const_source (

            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),

            .HI(one_unbuf),
            .LO(zero_unbuf)
    );

    assign zero = zero_unbuf;
    assign one = one_unbuf;

endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

// This module represents an unprogrammed set of GPIO pad default
// values that is configured with via programming on the chip top
// level.  This value is passed as a set of parameters (formerly
// part of gpio_control_block.v).

module gpio_defaults_block #(
    // Parameterized initial startup state of the pad.  The default
    // parameters if unspecified is for the pad to be a user input
    // with no pull-up or pull-down, so that it is disconnected
    // from the outside world.  See defs.h for configuration word
    // definitions.
    parameter GPIO_CONFIG_INIT = 13'h0402
) (

    inout VPWR,
    inout VGND,

    output [12:0] gpio_defaults
);
    wire [12:0] gpio_defaults_high;
    wire [12:0] gpio_defaults_low;

    // For the mask revision input, use an array of digital constant logic cells

    sky130_fd_sc_hd__conb_1 gpio_default_value [12:0] (

            .VPWR(VPWR),
            .VPB(VPWR),
            .VNB(VGND),
            .VGND(VGND),

            .HI(gpio_defaults_high),
            .LO(gpio_defaults_low)
    );

    genvar i;
    generate
        for (i = 0; i < 13; i = i+1) begin
    	    assign gpio_defaults[i] = (GPIO_CONFIG_INIT & (13'h0001 << i)) ?
			gpio_defaults_high[i] : gpio_defaults_low[i];
	end
    endgenerate

endmodule
`default_nettype wire
module gpio_logic_high(
 
         inout vccd1,
         inout vssd1,
  

   output wire gpio_logic1
);

 sky130_fd_sc_hd__conb_1 gpio_logic_high (

            .VPWR(vccd1),
            .VGND(vssd1),
            .VPB(vccd1),
            .VNB(vssd1),

            .HI(gpio_logic1),
            .LO()
    );

endmodule
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/* 
 *---------------------------------------------------------------------
 * A simple module that generates buffered high and low outputs
 * in the 1.8V domain.
 *---------------------------------------------------------------------
 */

module constant_block (
    
         inout vccd,
         inout vssd,
    

    output	 one,
    output	 zero
);

    wire	one_unbuf;
    wire	zero_unbuf;

    sky130_fd_sc_hd__conb_1 const_source (

            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),

            .HI(one_unbuf),
            .LO(zero_unbuf)
    );

    /* Buffer the constant outputs (could be synthesized) */
    /* NOTE:  Constant cell HI, LO outputs are connected to power	*/
    /* rails through an approximately 120 ohm resistor, which is not	*/
    /* enough to drive inputs in the I/O cells while ensuring ESD	*/
    /* requirements, without buffering.					*/

    sky130_fd_sc_hd__buf_16 const_one_buf (

            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),

            .A(one_unbuf),
            .X(one)
    );

    sky130_fd_sc_hd__buf_16 const_zero_buf (

            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),

            .A(zero_unbuf),
            .X(zero)
    );

endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// Module xres_buf is a level-shift buffer between the xres pad (used for
// digital reset) and the caravel chip core.  The xres pad output is in
// the 3.3V domain while the signal goes to the digital circuitry in the
// 1.8V domain.

module xres_buf (
	X    ,
	A    ,

	VPWR ,
	VGND ,
	LVPWR,
	LVGND,

);

output X    ;
input  A    ;

inout  VPWR ;
inout  VGND ;
inout  LVPWR;
inout  LVGND;


sky130_fd_sc_hvl__lsbufhv2lv_1 lvlshiftdown (

	.VPWR(VPWR),
	.VPB(VPWR),

	.LVPWR(LVPWR),

	.VNB(VGND),
	.VGND(VGND),

	.A(A),
	.X(X)
);

endmodule
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

// Spare logic block.  This block can be used for metal mask fixes to
// a design.  It is much larger and more comprehensive than the simple
// "macro_sparecell" in the HD library, and contains flops, taps, muxes,
// and diodes in addition to the inverters, NOR, NAND, and constant
// gates provided by macro_sparecell.

module spare_logic_block (
    
        inout vccd,
        inout vssd,
    

    output [26:0] spare_xz,	// Constant 0 outputs (and block inputs)
    output [3:0]  spare_xi,	// Inverter outputs
    output	  spare_xib,	// Big inverter output
    output [1:0]  spare_xna,	// NAND outputs
    output [1:0]  spare_xno,	// NOR outputs
    output [1:0]  spare_xmx,	// Mux outputs
    output [1:0]  spare_xfq,	// Flop noninverted output
    output [1:0]  spare_xfqn 	// Flop inverted output
);

    wire [3:0] spare_logic_nc;

    wire [26:0] spare_logic1;
    wire [26:0] spare_logic0;

    // Rename the logic0 outputs at the block pins.
    assign spare_xz = spare_logic0;

    sky130_fd_sc_hd__conb_1 spare_logic_const [26:0] (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
	
            .HI(spare_logic1),
            .LO(spare_logic0)
    );

    sky130_fd_sc_hd__inv_2 spare_logic_inv [3:0] (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
	
            .Y(spare_xi),
            .A(spare_logic0[3:0])
    );

    sky130_fd_sc_hd__inv_8 spare_logic_biginv (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
	
            .Y(spare_xib),
            .A(spare_logic0[4])
    );

    sky130_fd_sc_hd__nand2_2 spare_logic_nand [1:0] (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
	
            .Y(spare_xna),
            .A(spare_logic0[6:5]),
            .B(spare_logic0[8:7])
    );

    sky130_fd_sc_hd__nor2_2 spare_logic_nor [1:0] (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
	
            .Y(spare_xno),
            .A(spare_logic0[10:9]),
            .B(spare_logic0[12:11])
    );

    sky130_fd_sc_hd__mux2_2 spare_logic_mux [1:0] (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
	
            .X(spare_xmx),
            .A0(spare_logic0[14:13]),
            .A1(spare_logic0[16:15]),
            .S(spare_logic0[18:17])
    );

    sky130_fd_sc_hd__dfbbp_1 spare_logic_flop [1:0] (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
	
            .Q(spare_xfq),
            .Q_N(spare_xfqn),
            .D(spare_logic0[20:19]),
            .CLK(spare_logic0[22:21]),
            .SET_B(spare_logic0[24:23]),
            .RESET_B(spare_logic0[26:25])
    );

    sky130_fd_sc_hd__tapvpwrvgnd_1 spare_logic_tap [1:0] (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd)
	
    );

    sky130_fd_sc_hd__diode_2 spare_logic_diode [3:0] (
	
            .VPWR(vccd),
            .VGND(vssd),
            .VPB(vccd),
            .VNB(vssd),
	
	    .DIODE(spare_logic_nc)
    );
 
endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

//-----------------------------------------------------------
// Housekeeping interface for Caravel
//-----------------------------------------------------------
// Written by Tim Edwards
// efabless, inc. September 27, 2020
//-----------------------------------------------------------

//-----------------------------------------------------------
// This is a standalone slave SPI for the caravel chip that is
// intended to be independent of the picosoc and independent
// of all IP blocks except the power-on-reset.  This SPI has
// register outputs controlling the functions that critically
// affect operation of the picosoc and so cannot be accessed
// from the picosoc itself.  This includes the PLL enables,
// mode, and trim.  It also has a general reset for the picosoc,
// an IRQ input, a bypass for the entire crystal oscillator
// and PLL chain, the manufacturer and product IDs and product
// revision number.
//
// Updated and revised, 10/13/2021:
// This module now comprises what was previously split into
// the housekeeping SPI, the mprj_ctrl block (control over
// the GPIO), and sysctrl (redirection of certain internal
// signals to the GPIO);  and additionally manages the SPI
// flash signals and pass-through mode.  Essentially all
// aspects of the system related to the use and configuration
// of the GPIO has been shifted to this module.  This allows
// GPIO to be configured from either the management SoC
// through the wishbone interface, or externally through the
// SPI interface.  It allows essentially any processor to
// take the place of the PicoRV32 as long as that processor
// can access memory-mapped space via the wishbone bus.
//-----------------------------------------------------------

//------------------------------------------------------------
// Caravel defined registers (by SPI address):
// See:  doc/memory_map.txt
//------------------------------------------------------------

module housekeeping #(
    parameter GPIO_BASE_ADR = 32'h2600_0000,
    parameter SPI_BASE_ADR = 32'h2610_0000,
    parameter SYS_BASE_ADR = 32'h2620_0000,
    parameter IO_CTRL_BITS = 13
) (

    inout VPWR,
    inout VGND, 


    // Wishbone interface to management SoC
    input wb_clk_i,
    input wb_rstn_i,
    input [31:0] wb_adr_i,
    input [31:0] wb_dat_i,
    input [3:0] wb_sel_i,
    input wb_we_i,
    input wb_cyc_i,
    input wb_stb_i,
    output reg wb_ack_o,
    output reg [31:0] wb_dat_o,

    // Primary reset
    input porb,

    // Clocking control parameters
    output reg pll_ena,
    output reg pll_dco_ena,
    output reg [4:0] pll_div,
    output reg [2:0] pll_sel,
    output reg [2:0] pll90_sel,
    output reg [25:0] pll_trim,
    output reg pll_bypass,

    // Module enable status from SoC
    input  qspi_enabled,	// Flash SPI is in quad mode
    input  uart_enabled,	// UART is enabled
    input  spi_enabled,		// SPI master is enabled
    input  debug_mode,		// Debug mode enabled

    // UART interface to/from SoC
    input  ser_tx,
    output ser_rx,

    // SPI master interface to/from SoC
    output spi_sdi,
    input  spi_csb,
    input  spi_sck,
    input  spi_sdo,
    input  spi_sdoenb,

    // External (originating from SPI and pad) IRQ and reset
    output [2:0] irq,
    output reset,

    // GPIO serial loader programming interface
    output serial_clock,
    output serial_load,
    output serial_resetn,
    output serial_data_1,
    output serial_data_2,

    // GPIO data management (to padframe)---three-pin interface
    input  [(19 + 19)-1:0] mgmt_gpio_in,
    output [(19 + 19)-1:0] mgmt_gpio_out,
    output [(19 + 19)-1:0] mgmt_gpio_oeb,

    // Power control output (reserved for future use with LDOs)
    output reg [(2 + 2)-1:0] pwr_ctrl_out,

    // CPU trap state status (for system monitoring)
    input trap,

    // User clock (for system monitoring)
    input user_clock,

    // Mask revision/User project ID
    input [31:0] mask_rev_in,

    // SPI flash management (management SoC side)
    input spimemio_flash_csb,
    input spimemio_flash_clk,
    input spimemio_flash_io0_oeb,
    input spimemio_flash_io1_oeb,
    input spimemio_flash_io2_oeb,
    input spimemio_flash_io3_oeb,
    input spimemio_flash_io0_do,
    input spimemio_flash_io1_do,
    input spimemio_flash_io2_do,
    input spimemio_flash_io3_do,
    output spimemio_flash_io0_di,
    output spimemio_flash_io1_di,
    output spimemio_flash_io2_di,
    output spimemio_flash_io3_di,

    // Debug interface (routes to first GPIO) from management SoC
    output debug_in,
    input debug_out,
    input debug_oeb,

    // SPI flash management (padframe side)
    // (io2 and io3 are part of GPIO array, not dedicated pads)
    output pad_flash_csb,
    output pad_flash_csb_oeb,
    output pad_flash_clk,
    output pad_flash_clk_oeb,
    output pad_flash_io0_oeb,
    output pad_flash_io1_oeb,
    output pad_flash_io0_ieb,
    output pad_flash_io1_ieb,
    output pad_flash_io0_do,
    output pad_flash_io1_do,
    input pad_flash_io0_di,
    input pad_flash_io1_di,








    // System signal monitoring
    input  usr1_vcc_pwrgood,
    input  usr2_vcc_pwrgood,
    input  usr1_vdd_pwrgood,
    input  usr2_vdd_pwrgood
);

    localparam OEB = 1;		// Offset of output enable (bar) in shift register
    localparam INP_DIS = 3;	// Offset of input disable in shift register

    reg reset_reg;
    reg irq_spi;
    reg serial_bb_clock;
    reg serial_bb_load;
    reg serial_bb_resetn;
    reg serial_bb_data_1;
    reg serial_bb_data_2;
    reg serial_bb_enable;
    reg serial_xfer;
    reg hkspi_disable;







    reg clk1_output_dest;
    reg clk2_output_dest;
    reg trap_output_dest;
    reg irq_1_inputsrc;
    reg irq_2_inputsrc;

    reg [IO_CTRL_BITS-1:0] gpio_configure [(19 + 19)-1:0];
    reg [(19 + 19)-1:0] mgmt_gpio_data;

    /* mgmt_gpio_data_buf holds the lower bits during a back-door
     * write to GPIO data so that all 32 bits can update at once.
     */
    reg [23:0] mgmt_gpio_data_buf;


    wire [7:0] odata;
    wire [7:0] idata;
    wire [7:0] iaddr;

    wire rdstb;
    wire wrstb;
    wire pass_thru_mgmt;		// Mode detected by housekeeping_spi
    wire pass_thru_mgmt_delay;
    wire pass_thru_user;		// Mode detected by housekeeping_spi
    wire pass_thru_user_delay;
    wire pass_thru_mgmt_reset;
    wire pass_thru_user_reset;
    wire sdo;
    wire sdo_enb;

    wire [7:0]	caddr;	// Combination of SPI address and back door address
    wire [7:0]	cdata;	// Combination of SPI data and back door data
    wire	cwstb;	// Combination of SPI write strobe and back door write strobe
    wire	csclk;	// Combination of SPI SCK and back door access trigger


// Output clock signals buffer wires
wire mgmt_gpio_out_9_prebuff, mgmt_gpio_out_14_prebuff, mgmt_gpio_out_15_prebuff, pad_flash_clk_prebuff;






    // Pass-through mode handling.  Signals may only be applied when the
    // core processor is in reset.

    assign reset = (pass_thru_mgmt_reset) ? 1'b1 : reset_reg;

	// Invert wb_rstn_i
	wire wb_rst_i;
	assign wb_rst_i = ~wb_rstn_i;
	
    // Pass-through mode.  Housekeeping SPI signals get inserted
    // between the management SoC and the flash SPI I/O.

    assign pad_flash_csb = (pass_thru_mgmt_delay) ? mgmt_gpio_in[3] : spimemio_flash_csb;
    assign pad_flash_csb_oeb = (pass_thru_mgmt_delay) ? 1'b0 : (~porb ? 1'b1 : 1'b0);
    assign pad_flash_clk_prebuff = (pass_thru_mgmt) ? mgmt_gpio_in[4] : spimemio_flash_clk;
    assign pad_flash_clk_oeb = (pass_thru_mgmt) ? 1'b0 : (~porb ? 1'b1 : 1'b0);
    assign pad_flash_io0_oeb = (pass_thru_mgmt_delay) ? 1'b0 : spimemio_flash_io0_oeb;
    assign pad_flash_io1_oeb = (pass_thru_mgmt) ? 1'b1 : spimemio_flash_io1_oeb;
    assign pad_flash_io0_ieb = (pass_thru_mgmt_delay) ? 1'b1 : ~spimemio_flash_io0_oeb;
    assign pad_flash_io1_ieb = (pass_thru_mgmt) ? 1'b0 : ~spimemio_flash_io1_oeb;
    assign pad_flash_io0_do = (pass_thru_mgmt_delay) ? mgmt_gpio_in[2] : spimemio_flash_io0_do;
    assign pad_flash_io1_do = spimemio_flash_io1_do;
    assign spimemio_flash_io0_di = (pass_thru_mgmt_delay) ? 1'b0 : pad_flash_io0_di;
    assign spimemio_flash_io1_di = (pass_thru_mgmt) ? 1'b0 : pad_flash_io1_di;

(* keep *) sky130_fd_sc_hd__clkbuf_8 pad_flashh_clk_buff_inst (

        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPWR),
        .VNB(VGND),

	.A(pad_flash_clk_prebuff),
    .X(pad_flash_clk));

    wire [11:0] mfgr_id;
    wire [7:0]  prod_id;
    wire [31:0] mask_rev;

    reg serial_busy;

    // Wishbone bus "back door" to SPI registers.  This section of code
    // (1) Maps SPI byte addresses to memory map 32-bit addresses
    // (2) Applies signals to the housekeeping SPI to mux in the SPI address,
    //	   clock, and write strobe.  This is done carefully and slowly to
    //	   avoid glitching on the SCK line and to avoid forcing the
    //	   housekeeping module to keep up with the core clock timing.

    wire      	sys_select;	// System monitoring memory map address selected
    wire      	gpio_select;	// GPIO configuration memory map address selected
    wire      	spi_select;	// SPI back door memory map address selected

    // Wishbone Back Door.  This is a simple interface making use of the
    // housekeeping SPI protocol.  The housekeeping SPI uses byte-wide
    // data, so this interface will stall the processor by holding wb_ack_o
    // low until all bytes have been transferred between the processor and
    // housekeeping SPI.

    reg [3:0] 	wbbd_state;
    reg [7:0] 	wbbd_addr;	/* SPI address translated from WB */
    reg [7:0] 	wbbd_data;	/* SPI data translated from WB */
    reg  	wbbd_sck;	/* wishbone access trigger (back-door clock) */
    reg  	wbbd_write;	/* wishbone write trigger (back-door strobe) */
    reg		wbbd_busy;	/* Raised during a wishbone read or write */

    // This defines a state machine that accesses the SPI registers through
    // the back door wishbone interface.  The process is relatively slow
    // since the SPI data are byte-wide, so four individual accesses are
    // made to read 4 bytes from the SPI to fill data on the wishbone bus
    // before sending ACK and letting the processor continue.

    
    
    
    
    
    
    
    
    
    
    

    assign sys_select = (wb_adr_i[31:8] == SYS_BASE_ADR[31:8]);
    assign gpio_select = (wb_adr_i[31:8] == GPIO_BASE_ADR[31:8]);
    assign spi_select = (wb_adr_i[31:8] == SPI_BASE_ADR[31:8]);

    /* Register bit to SPI address mapping */

    function [7:0] fdata(input [7:0] address);
	begin
	case (address)
	    /* Housekeeping SPI Protocol */
	    8'h00 : fdata = 8'h00;			// SPI status (fixed) 

	    /* Status and Identification */
	    8'h01 : fdata = {4'h0, mfgr_id[11:8]};	// Manufacturer ID (fixed)
	    8'h02 : fdata = mfgr_id[7:0];		// Manufacturer ID (fixed)
	    8'h03 : fdata = prod_id;			// Product ID (fixed)
	    8'h04 : fdata = mask_rev[31:24];		// Mask rev (via programmed)
	    8'h05 : fdata = mask_rev[23:16];		// Mask rev (via programmed)
	    8'h06 : fdata = mask_rev[15:8];		// Mask rev (via programmed)
	    8'h07 : fdata = mask_rev[7:0];		// Mask rev (via programmed)

	    /* Clocking control */
	    8'h08 : fdata = {6'b000000, pll_dco_ena, pll_ena};
	    8'h09 : fdata = {7'b0000000, pll_bypass};
	    8'h0a : fdata = {7'b0000000, irq_spi};
	    8'h0b : fdata = {7'b0000000, reset};
	    8'h0c : fdata = {7'b0000000, trap};		// CPU trap state
	    8'h0d : fdata = pll_trim[7:0];
	    8'h0e : fdata = pll_trim[15:8];
	    8'h0f : fdata = pll_trim[23:16];
	    8'h10 : fdata = {6'b000000, pll_trim[25:24]};
	    8'h11 : fdata = {2'b00, pll90_sel, pll_sel};
	    8'h12 : fdata = {3'b000, pll_div};

	    // GPIO Control (bit bang and automatic)
	    // NOTE: "serial_busy" is the read-back signal occupying the same
	    // address/bit as "serial_xfer".
	    8'h13 : fdata = {1'b0, serial_data_2, serial_data_1, serial_bb_clock,
				serial_bb_load, serial_bb_resetn, serial_bb_enable,
				serial_busy};











	    /* System monitoring */
	    8'h1a : fdata = {4'b0000, usr1_vcc_pwrgood, usr2_vcc_pwrgood,
				usr1_vdd_pwrgood, usr2_vdd_pwrgood};
	    8'h1b : fdata = {5'b00000, clk1_output_dest, clk2_output_dest,
				trap_output_dest};
	    8'h1c : fdata = {6'b000000, irq_2_inputsrc, irq_1_inputsrc};

	    /* GPIO Configuration */
	    8'h1d : fdata = {3'b000, gpio_configure[0][12:8]};
	    8'h1e : fdata = gpio_configure[0][7:0];
	    8'h1f : fdata = {3'b000, gpio_configure[1][12:8]};
	    8'h20 : fdata = gpio_configure[1][7:0];
	    8'h21 : fdata = {3'b000, gpio_configure[2][12:8]};
	    8'h22 : fdata = gpio_configure[2][7:0];
	    8'h23 : fdata = {3'b000, gpio_configure[3][12:8]};
	    8'h24 : fdata = gpio_configure[3][7:0];
	    8'h25 : fdata = {3'b000, gpio_configure[4][12:8]};
	    8'h26 : fdata = gpio_configure[4][7:0];
	    8'h27 : fdata = {3'b000, gpio_configure[5][12:8]};
	    8'h28 : fdata = gpio_configure[5][7:0];
	    8'h29 : fdata = {3'b000, gpio_configure[6][12:8]};
	    8'h2a : fdata = gpio_configure[6][7:0];
	    8'h2b : fdata = {3'b000, gpio_configure[7][12:8]};
	    8'h2c : fdata = gpio_configure[7][7:0];
	    8'h2d : fdata = {3'b000, gpio_configure[8][12:8]};
	    8'h2e : fdata = gpio_configure[8][7:0];
	    8'h2f : fdata = {3'b000, gpio_configure[9][12:8]};
	    8'h30 : fdata = gpio_configure[9][7:0];
	    8'h31 : fdata = {3'b000, gpio_configure[10][12:8]};
	    8'h32 : fdata = gpio_configure[10][7:0];
	    8'h33 : fdata = {3'b000, gpio_configure[11][12:8]};
	    8'h34 : fdata = gpio_configure[11][7:0];
	    8'h35 : fdata = {3'b000, gpio_configure[12][12:8]};
	    8'h36 : fdata = gpio_configure[12][7:0];
	    8'h37 : fdata = {3'b000, gpio_configure[13][12:8]};
	    8'h38 : fdata = gpio_configure[13][7:0];
	    8'h39 : fdata = {3'b000, gpio_configure[14][12:8]};
	    8'h3a : fdata = gpio_configure[14][7:0];
	    8'h3b : fdata = {3'b000, gpio_configure[15][12:8]};
	    8'h3c : fdata = gpio_configure[15][7:0];
	    8'h3d : fdata = {3'b000, gpio_configure[16][12:8]};
	    8'h3e : fdata = gpio_configure[16][7:0];
	    8'h3f : fdata = {3'b000, gpio_configure[17][12:8]};
	    8'h40 : fdata = gpio_configure[17][7:0];
	    8'h41 : fdata = {3'b000, gpio_configure[18][12:8]};
	    8'h42 : fdata = gpio_configure[18][7:0];
	    8'h43 : fdata = {3'b000, gpio_configure[19][12:8]};
	    8'h44 : fdata = gpio_configure[19][7:0];
	    8'h45 : fdata = {3'b000, gpio_configure[20][12:8]};
	    8'h46 : fdata = gpio_configure[20][7:0];
	    8'h47 : fdata = {3'b000, gpio_configure[21][12:8]};
	    8'h48 : fdata = gpio_configure[21][7:0];
	    8'h49 : fdata = {3'b000, gpio_configure[22][12:8]};
	    8'h4a : fdata = gpio_configure[22][7:0];
	    8'h4b : fdata = {3'b000, gpio_configure[23][12:8]};
	    8'h4c : fdata = gpio_configure[23][7:0];
	    8'h4d : fdata = {3'b000, gpio_configure[24][12:8]};
	    8'h4e : fdata = gpio_configure[24][7:0];
	    8'h4f : fdata = {3'b000, gpio_configure[25][12:8]};
	    8'h50 : fdata = gpio_configure[25][7:0];
	    8'h51 : fdata = {3'b000, gpio_configure[26][12:8]};
	    8'h52 : fdata = gpio_configure[26][7:0];
	    8'h53 : fdata = {3'b000, gpio_configure[27][12:8]};
	    8'h54 : fdata = gpio_configure[27][7:0];
	    8'h55 : fdata = {3'b000, gpio_configure[28][12:8]};
	    8'h56 : fdata = gpio_configure[28][7:0];
	    8'h57 : fdata = {3'b000, gpio_configure[29][12:8]};
	    8'h58 : fdata = gpio_configure[29][7:0];
	    8'h59 : fdata = {3'b000, gpio_configure[30][12:8]};
	    8'h5a : fdata = gpio_configure[30][7:0];
	    8'h5b : fdata = {3'b000, gpio_configure[31][12:8]};
	    8'h5c : fdata = gpio_configure[31][7:0];
	    8'h5d : fdata = {3'b000, gpio_configure[32][12:8]};
	    8'h5e : fdata = gpio_configure[32][7:0];
	    8'h5f : fdata = {3'b000, gpio_configure[33][12:8]};
	    8'h60 : fdata = gpio_configure[33][7:0];
	    8'h61 : fdata = {3'b000, gpio_configure[34][12:8]};
	    8'h62 : fdata = gpio_configure[34][7:0];
	    8'h63 : fdata = {3'b000, gpio_configure[35][12:8]};
	    8'h64 : fdata = gpio_configure[35][7:0];
	    8'h65 : fdata = {3'b000, gpio_configure[36][12:8]};
	    8'h66 : fdata = gpio_configure[36][7:0];
	    8'h67 : fdata = {3'b000, gpio_configure[37][12:8]};
	    8'h68 : fdata = gpio_configure[37][7:0];

	    // GPIO Data
	    8'h69 : fdata = {2'b00, mgmt_gpio_in[(19 + 19)-1:32]};
	    8'h6a : fdata = mgmt_gpio_in[31:24];
	    8'h6b : fdata = mgmt_gpio_in[23:16];
	    8'h6c : fdata = mgmt_gpio_in[15:8];
	    8'h6d : fdata = mgmt_gpio_in[7:0];

	    // Power Control (reserved)
	    8'h6e : fdata = {4'b0000, pwr_ctrl_out};

	    // Housekeeping SPI system disable
	    8'h6f : fdata = {7'b0000000, hkspi_disable};

	    default: fdata = 8'h00;
	endcase
	end
    endfunction

    /* Memory map address to SPI address translation for back door access */
    /* (see doc/memory_map.txt)						  */

    wire [11:0] gpio_adr = GPIO_BASE_ADR[23:12];
    wire [11:0] sys_adr = SYS_BASE_ADR[23:12];
    wire [11:0] spi_adr = SPI_BASE_ADR[23:12];

    function [7:0] spiaddr(input [31:0] wbaddress);
	begin
	/* Address taken from lower 8 bits and upper 4 bits of the 32-bit */
	/* wishbone address.						  */
	case ({wbaddress[23:20], wbaddress[7:0]})
	    spi_adr  | 12'h000 : spiaddr = 8'h00;	// SPI status (reserved)
	    spi_adr  | 12'h004 : spiaddr = 8'h03;	// product ID
	    spi_adr  | 12'h005 : spiaddr = 8'h02;	// Manufacturer ID (low)
	    spi_adr  | 12'h006 : spiaddr = 8'h01;	// Manufacturer ID (high)
	    spi_adr  | 12'h008 : spiaddr = 8'h07;	// User project ID (low)
	    spi_adr  | 12'h009 : spiaddr = 8'h06;	// User project ID .
	    spi_adr  | 12'h00a : spiaddr = 8'h05;	// User project ID .
	    spi_adr  | 12'h00b : spiaddr = 8'h04;	// User project ID (high)

	    spi_adr  | 12'h00c : spiaddr = 8'h08;	// PLL enables
	    spi_adr  | 12'h010 : spiaddr = 8'h09;	// PLL bypass
	    spi_adr  | 12'h014 : spiaddr = 8'h0a;	// IRQ
	    spi_adr  | 12'h018 : spiaddr = 8'h0b;	// Reset
	    spi_adr  | 12'h028 : spiaddr = 8'h0c;	// CPU trap state
	    spi_adr  | 12'h01f : spiaddr = 8'h10;	// PLL trim
	    spi_adr  | 12'h01e : spiaddr = 8'h0f;	// PLL trim
	    spi_adr  | 12'h01d : spiaddr = 8'h0e;	// PLL trim
	    spi_adr  | 12'h01c : spiaddr = 8'h0d;	// PLL trim
	    spi_adr  | 12'h020 : spiaddr = 8'h11;	// PLL source
	    spi_adr  | 12'h024 : spiaddr = 8'h12;	// PLL divider

	    spi_adr  | 12'h02c : spiaddr = 8'h19;	// SRAM read-only data
	    spi_adr  | 12'h02d : spiaddr = 8'h18;	// SRAM read-only data
	    spi_adr  | 12'h02e : spiaddr = 8'h17;	// SRAM read-only data
	    spi_adr  | 12'h02f : spiaddr = 8'h16;	// SRAM read-only data
	    spi_adr  | 12'h030 : spiaddr = 8'h15;	// SRAM read-only address
	    spi_adr  | 12'h034 : spiaddr = 8'h14;	// SRAM read-only control

	    gpio_adr | 12'h000 : spiaddr = 8'h13;	// GPIO control

	    sys_adr  | 12'h000 : spiaddr = 8'h1a;	// Power monitor
	    sys_adr  | 12'h004 : spiaddr = 8'h1b;	// Output redirect
	    sys_adr  | 12'h00c : spiaddr = 8'h1c;	// Input redirect

	    gpio_adr | 12'h025 : spiaddr = 8'h1d;	// GPIO configuration
	    gpio_adr | 12'h024 : spiaddr = 8'h1e;
	    gpio_adr | 12'h029 : spiaddr = 8'h1f;
	    gpio_adr | 12'h028 : spiaddr = 8'h20;
	    gpio_adr | 12'h02d : spiaddr = 8'h21;
	    gpio_adr | 12'h02c : spiaddr = 8'h22;
	    gpio_adr | 12'h031 : spiaddr = 8'h23;
	    gpio_adr | 12'h030 : spiaddr = 8'h24;
	    gpio_adr | 12'h035 : spiaddr = 8'h25;
	    gpio_adr | 12'h034 : spiaddr = 8'h26;
	    gpio_adr | 12'h039 : spiaddr = 8'h27;
	    gpio_adr | 12'h038 : spiaddr = 8'h28;
	    gpio_adr | 12'h03d : spiaddr = 8'h29;
	    gpio_adr | 12'h03c : spiaddr = 8'h2a;
	    gpio_adr | 12'h041 : spiaddr = 8'h2b;
	    gpio_adr | 12'h040 : spiaddr = 8'h2c;
	    gpio_adr | 12'h045 : spiaddr = 8'h2d;
	    gpio_adr | 12'h044 : spiaddr = 8'h2e;
	    gpio_adr | 12'h049 : spiaddr = 8'h2f;
	    gpio_adr | 12'h048 : spiaddr = 8'h30;
	    gpio_adr | 12'h04d : spiaddr = 8'h31;
	    gpio_adr | 12'h04c : spiaddr = 8'h32;
	    gpio_adr | 12'h051 : spiaddr = 8'h33;
	    gpio_adr | 12'h050 : spiaddr = 8'h34;
	    gpio_adr | 12'h055 : spiaddr = 8'h35;
	    gpio_adr | 12'h054 : spiaddr = 8'h36;
	    gpio_adr | 12'h059 : spiaddr = 8'h37;
	    gpio_adr | 12'h058 : spiaddr = 8'h38;
	    gpio_adr | 12'h05d : spiaddr = 8'h39;
	    gpio_adr | 12'h05c : spiaddr = 8'h3a;
	    gpio_adr | 12'h061 : spiaddr = 8'h3b;
	    gpio_adr | 12'h060 : spiaddr = 8'h3c;
	    gpio_adr | 12'h065 : spiaddr = 8'h3d;
	    gpio_adr | 12'h064 : spiaddr = 8'h3e;
	    gpio_adr | 12'h069 : spiaddr = 8'h3f;
	    gpio_adr | 12'h068 : spiaddr = 8'h40;
	    gpio_adr | 12'h06d : spiaddr = 8'h41;
	    gpio_adr | 12'h06c : spiaddr = 8'h42;
	    gpio_adr | 12'h071 : spiaddr = 8'h43;
	    gpio_adr | 12'h070 : spiaddr = 8'h44;
	    gpio_adr | 12'h075 : spiaddr = 8'h45;
	    gpio_adr | 12'h074 : spiaddr = 8'h46;
	    gpio_adr | 12'h079 : spiaddr = 8'h47;
	    gpio_adr | 12'h078 : spiaddr = 8'h48;
	    gpio_adr | 12'h07d : spiaddr = 8'h49;
	    gpio_adr | 12'h07c : spiaddr = 8'h4a;
	    gpio_adr | 12'h081 : spiaddr = 8'h4b;
	    gpio_adr | 12'h080 : spiaddr = 8'h4c;
	    gpio_adr | 12'h085 : spiaddr = 8'h4d;
	    gpio_adr | 12'h084 : spiaddr = 8'h4e;
	    gpio_adr | 12'h089 : spiaddr = 8'h4f;
	    gpio_adr | 12'h088 : spiaddr = 8'h50;
	    gpio_adr | 12'h08d : spiaddr = 8'h51;
	    gpio_adr | 12'h08c : spiaddr = 8'h52;
	    gpio_adr | 12'h091 : spiaddr = 8'h53;
	    gpio_adr | 12'h090 : spiaddr = 8'h54;
	    gpio_adr | 12'h095 : spiaddr = 8'h55;
	    gpio_adr | 12'h094 : spiaddr = 8'h56;
	    gpio_adr | 12'h099 : spiaddr = 8'h57;
	    gpio_adr | 12'h098 : spiaddr = 8'h58;
	    gpio_adr | 12'h09d : spiaddr = 8'h59;
	    gpio_adr | 12'h09c : spiaddr = 8'h5a;
	    gpio_adr | 12'h0a1 : spiaddr = 8'h5b;
	    gpio_adr | 12'h0a0 : spiaddr = 8'h5c;
	    gpio_adr | 12'h0a5 : spiaddr = 8'h5d;
	    gpio_adr | 12'h0a4 : spiaddr = 8'h5e;
	    gpio_adr | 12'h0a9 : spiaddr = 8'h5f;
	    gpio_adr | 12'h0a8 : spiaddr = 8'h60;
	    gpio_adr | 12'h0ad : spiaddr = 8'h61;
	    gpio_adr | 12'h0ac : spiaddr = 8'h62;
	    gpio_adr | 12'h0b1 : spiaddr = 8'h63;
	    gpio_adr | 12'h0b0 : spiaddr = 8'h64;
	    gpio_adr | 12'h0b5 : spiaddr = 8'h65;
	    gpio_adr | 12'h0b4 : spiaddr = 8'h66;
	    gpio_adr | 12'h0b9 : spiaddr = 8'h67;
	    gpio_adr | 12'h0b8 : spiaddr = 8'h68;

	    gpio_adr | 12'h010 : spiaddr = 8'h69;	// GPIO data (h)

	    gpio_adr | 12'h00f : spiaddr = 8'h6a;	// GPIO data (l)
	    gpio_adr | 12'h00e : spiaddr = 8'h6b;	// GPIO data (l)
	    gpio_adr | 12'h00d : spiaddr = 8'h6c;	// GPIO data (l)
	    gpio_adr | 12'h00c : spiaddr = 8'h6d;	// GPIO data (l)

	    gpio_adr | 12'h004 : spiaddr = 8'h6e;	// Power control

	    sys_adr  | 12'h010 : spiaddr = 8'h6f;	// Housekeeping SPI disable

	    default : spiaddr = 8'h00;
	endcase
	end
    endfunction
	
    // SPI is considered active when the GPIO for CSB is set to input and
    // CSB is low.  SPI is considered "busy" when rdstb or wrstb are high,
    // indicating that the SPI will read or write a byte on the next SCK
    // transition.

    wire spi_is_enabled = (~gpio_configure[3][INP_DIS]) & (~hkspi_disable);
    wire spi_is_active = spi_is_enabled && (mgmt_gpio_in[3] == 1'b0);
    wire spi_is_busy = spi_is_active && (rdstb || wrstb);

    /* Wishbone back-door state machine and address translation */

    always @(posedge wb_clk_i or posedge wb_rst_i) begin
	if (wb_rst_i) begin
	    wbbd_sck <= 1'b0;
	    wbbd_write <= 1'b0;
	    wbbd_addr <= 8'd0;
	    wbbd_data <= 8'd0;
	    wbbd_busy <= 1'b0;
	    wb_ack_o <= 1'b0;
	    wbbd_state <= 4'h0;
	end else begin
	    case (wbbd_state)
		4'h0: begin
		    wbbd_sck <= 1'b0;
		    wbbd_busy <= 1'b0;
		    if ((sys_select | gpio_select | spi_select) &&
	    	    		 wb_cyc_i && wb_stb_i) begin
			wb_ack_o <= 1'b0;
			wbbd_state <= 4'h1;
		    end
		end
		4'h1: begin
		    wbbd_sck <= 1'b0;
		    wbbd_addr <= spiaddr(wb_adr_i);
		    if (wb_sel_i[0] & wb_we_i) begin
		    	wbbd_data <= wb_dat_i[7:0];
		    end
		    wbbd_write <= wb_sel_i[0] & wb_we_i;
		    wbbd_busy <= 1'b1;

		    // If the SPI is being accessed and about to read or
		    // write a byte, then stall until the SPI is ready.
		    if (!spi_is_busy) begin
		        wbbd_state <= 4'h2;
		    end
		end
		4'h2: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_dat_o[7:0] <= odata;
		    wbbd_state <= 4'h3;
		end
		4'h3: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b0;
		    wbbd_addr <= spiaddr(wb_adr_i + 1);
		    if (wb_sel_i[1] & wb_we_i) begin
		    	wbbd_data <= wb_dat_i[15:8];
		    end
		    wbbd_write <= wb_sel_i[1] & wb_we_i;
		    if (!spi_is_busy) begin
		        wbbd_state <= 4'h4;
		    end
		end
		4'h4: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_dat_o[15:8] <= odata;
		    wbbd_state <= 4'h5;
		end
		4'h5: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b0;
		    wbbd_addr <= spiaddr(wb_adr_i + 2);
		    if (wb_sel_i[2] & wb_we_i) begin
		    	wbbd_data <= wb_dat_i[23:16];
		    end
		    wbbd_write <= wb_sel_i[2] & wb_we_i;
		    if (!spi_is_busy) begin
		        wbbd_state <= 4'h6;
		    end
		end
		4'h6: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_dat_o[23:16] <= odata;
		    wbbd_state <= 4'h7;
		end
		4'h7: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b0;
		    wbbd_addr <= spiaddr(wb_adr_i + 3);
		    if (wb_sel_i[3] & wb_we_i) begin
		    	wbbd_data <= wb_dat_i[31:24];
		    end
		    wbbd_write <= wb_sel_i[3] & wb_we_i;
		    if (!spi_is_busy) begin
		        wbbd_state <= 4'h8;
		    end
		end
		4'h8: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_dat_o[31:24] <= odata;
		    wb_ack_o <= 1'b1;	// Release hold on wishbone bus
		    wbbd_state <= 4'h9;
		end
		4'h9: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b0;
		    wb_ack_o <= 1'b0;	// Reset for next access
		    wbbd_write <= 1'b0;
		    wbbd_state <= 4'ha;
		end
		4'ha: begin
		    wbbd_busy <= 1'b1;
		    wbbd_sck <= 1'b1;
		    wb_ack_o <= 1'b0;
		    wbbd_write <= 1'b0;
		    wbbd_state <= 4'h0;
		end
	    endcase
	end
    end

    // Instantiate the SPI interface protocol module

    housekeeping_spi hkspi (
	.reset(~porb),
    	.SCK(mgmt_gpio_in[4]),
    	.SDI(mgmt_gpio_in[2]),
    	.CSB((spi_is_enabled) ? mgmt_gpio_in[3] : 1'b1),
    	.SDO(sdo),
    	.sdoenb(sdo_enb),
    	.idata(odata),
    	.odata(idata),
    	.oaddr(iaddr),
    	.rdstb(rdstb),
    	.wrstb(wrstb),
    	.pass_thru_mgmt(pass_thru_mgmt),
    	.pass_thru_mgmt_delay(pass_thru_mgmt_delay),
    	.pass_thru_user(pass_thru_user),
    	.pass_thru_user_delay(pass_thru_user_delay),
    	.pass_thru_mgmt_reset(pass_thru_mgmt_reset),
    	.pass_thru_user_reset(pass_thru_user_reset)
    );



    // GPIO data handling to and from the management SoC

    assign mgmt_gpio_out[37] = (qspi_enabled) ? spimemio_flash_io3_do :
		mgmt_gpio_data[37];
    assign mgmt_gpio_out[36] = (qspi_enabled) ? spimemio_flash_io2_do :
		mgmt_gpio_data[36];

    assign mgmt_gpio_oeb[37] = (qspi_enabled) ? spimemio_flash_io3_oeb :
		~gpio_configure[37][INP_DIS];
    assign mgmt_gpio_oeb[36] = (qspi_enabled) ? spimemio_flash_io2_oeb :
		~gpio_configure[36][INP_DIS];
    assign mgmt_gpio_oeb[35] = (spi_enabled) ? spi_sdoenb :
		~gpio_configure[35][INP_DIS];

    // NOTE:  Ignored by spimemio module when QSPI disabled, so they do not
    // need any exception when qspi_enabled == 1.
    assign spimemio_flash_io3_di = mgmt_gpio_in[37];
    assign spimemio_flash_io2_di = mgmt_gpio_in[36];

    // SPI master is assigned to the other 4 bits of the data high word.
    assign mgmt_gpio_out[32] = (spi_enabled) ? spi_sck : mgmt_gpio_data[32];
    assign mgmt_gpio_out[33] = (spi_enabled) ? spi_csb : mgmt_gpio_data[33];
    assign mgmt_gpio_out[34] = mgmt_gpio_data[34];
    assign mgmt_gpio_out[35] = (spi_enabled) ? spi_sdo : mgmt_gpio_data[35];

    assign mgmt_gpio_out[31:16] = mgmt_gpio_data[31:16];
    assign mgmt_gpio_out[12:11] = mgmt_gpio_data[12:11];

    assign mgmt_gpio_out[10] = (pass_thru_user_delay) ? mgmt_gpio_in[2]
			: mgmt_gpio_data[10];
    assign mgmt_gpio_out_9_prebuff = (pass_thru_user) ? mgmt_gpio_in[4]
			: mgmt_gpio_data[9];

(* keep *) sky130_fd_sc_hd__clkbuf_8 mgmt_gpio_9_buff_inst (

        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPWR),
        .VNB(VGND),

	.A(mgmt_gpio_out_9_prebuff),
    .X(mgmt_gpio_out[9]));

    assign mgmt_gpio_out[8] = (pass_thru_user_delay) ? mgmt_gpio_in[3]
			: mgmt_gpio_data[8];

    assign mgmt_gpio_out[7] = mgmt_gpio_data[7];
    assign mgmt_gpio_out[6] = (uart_enabled) ? ser_tx : mgmt_gpio_data[6];
    assign mgmt_gpio_out[5:2] = mgmt_gpio_data[5:2];

    // In pass-through modes, route SDO from the respective flash (user or
    // management SoC) to the dedicated SDO pin (GPIO[1])

    assign mgmt_gpio_out[1] = (pass_thru_mgmt) ? pad_flash_io1_di :
		 (pass_thru_user) ? mgmt_gpio_in[11] :
		 (spi_is_active) ? sdo : mgmt_gpio_data[1];
    assign mgmt_gpio_out[0] = (debug_mode) ? debug_out : mgmt_gpio_data[0];

    assign mgmt_gpio_oeb[1] = (spi_is_active) ? sdo_enb : ~gpio_configure[1][INP_DIS];
    assign mgmt_gpio_oeb[0] = (debug_mode) ? debug_oeb : ~gpio_configure[0][INP_DIS];

    assign ser_rx = (uart_enabled) ? mgmt_gpio_in[5] : 1'b0;
    assign spi_sdi = (spi_enabled) ? mgmt_gpio_in[34] : 1'b0;
    assign debug_in = (debug_mode) ? mgmt_gpio_in[0] : 1'b0;

    genvar i;

    /* These are disconnected, but apply a meaningful signal anyway */
    generate
	for (i = 2; i < (19 + 19)-3; i = i + 1) begin
	    assign mgmt_gpio_oeb[i] = ~gpio_configure[i][INP_DIS];
	end
    endgenerate

    // System monitoring.  Multiplex the clock and trap
    // signals to the associated pad, and multiplex the irq signals
    // from the associated pad, when the redirection is enabled.  Note
    // that the redirection is upstream of the user/managment multiplexing,
    // so the pad being under control of the user area takes precedence
    // over the system monitoring function.

    assign mgmt_gpio_out_15_prebuff = (clk2_output_dest == 1'b1) ? user_clock
		: mgmt_gpio_data[15];

(* keep *) sky130_fd_sc_hd__clkbuf_8 mgmt_gpio_15_buff_inst (

        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPWR),
        .VNB(VGND),

	.A(mgmt_gpio_out_15_prebuff),
    .X(mgmt_gpio_out[15]));

    assign mgmt_gpio_out_14_prebuff = (clk1_output_dest == 1'b1) ? wb_clk_i
		: mgmt_gpio_data[14];

(* keep *) sky130_fd_sc_hd__clkbuf_8 mgmt_gpio_14_buff_inst (

        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPWR),
        .VNB(VGND),

	.A(mgmt_gpio_out_14_prebuff),
    .X(mgmt_gpio_out[14]));

    assign mgmt_gpio_out[13] = (trap_output_dest == 1'b1) ? trap
		: mgmt_gpio_data[13];

    assign irq[0] = irq_spi;
    assign irq[1] = (irq_1_inputsrc == 1'b1) ? mgmt_gpio_in[7] : 1'b0;
    assign irq[2] = (irq_2_inputsrc == 1'b1) ? mgmt_gpio_in[12] : 1'b0;

    // GPIO serial loader and GPIO management control






    reg [3:0]	xfer_count;
    reg [4:0]	pad_count_1;
    reg [5:0]	pad_count_2;
    reg [1:0]	xfer_state;

    reg serial_clock_pre;
    reg serial_resetn_pre;
    reg serial_load_pre;
    reg [IO_CTRL_BITS-1:0] serial_data_staging_1;
    reg [IO_CTRL_BITS-1:0] serial_data_staging_2;

    assign serial_clock = (serial_bb_enable == 1'b1) ?
			serial_bb_clock : serial_clock_pre;
    assign serial_resetn = (serial_bb_enable == 1'b1) ?
			serial_bb_resetn : serial_resetn_pre;
    assign serial_load = (serial_bb_enable == 1'b1) ?
			serial_bb_load : serial_load_pre;

    assign serial_data_1 = (serial_bb_enable == 1'b1) ?
			serial_bb_data_1 : serial_data_staging_1[IO_CTRL_BITS-1];
    assign serial_data_2 = (serial_bb_enable == 1'b1) ?
			serial_bb_data_2 : serial_data_staging_2[IO_CTRL_BITS-1];

    always @(posedge wb_clk_i or negedge porb) begin
	if (porb == 1'b0) begin
	    xfer_state <= 2'b00;
	    xfer_count <= 4'd0;
            /* NOTE:  This assumes that MPRJ_IO_PADS_1 and MPRJ_IO_PADS_2 are
             * equal, because they get clocked the same number of cycles by
             * the same clock signal.  pad_count_2 gates the count for both.
             */
	    pad_count_1 <= 19 - 1;
	    pad_count_2 <= 19;
	    serial_resetn_pre <= 1'b0;
	    serial_clock_pre <= 1'b0;
	    serial_load_pre <= 1'b0;
	    serial_data_staging_1 <= 0;
	    serial_data_staging_2 <= 0;
	    serial_busy <= 1'b0;

	end else begin

            serial_resetn_pre <= 1'b1;
	    case (xfer_state)
		2'b00: begin
		    pad_count_1 <= 19 - 1;
                    pad_count_2 <= 19;
                    serial_clock_pre <= 1'b0;
                    serial_load_pre <= 1'b0;
                    if (serial_xfer == 1'b1) begin
                        xfer_state <= 2'b01;
	    	    	serial_busy <= 1'b1;
                    end else begin
	    	    	serial_busy <= 1'b0;
		    end
		end
		2'b01: begin
                    serial_clock_pre <= 1'b0;
                    serial_load_pre <= 1'b0;
                    xfer_count <= 6'd0;
                    pad_count_1 <= pad_count_1 - 1;
                    pad_count_2 <= pad_count_2 + 1;
                    xfer_state <= 2'b10;
                    serial_data_staging_1 <= gpio_configure[pad_count_1];
                    serial_data_staging_2 <= gpio_configure[pad_count_2];
		end
		2'b10: begin
                    serial_clock_pre <= ~serial_clock;
                    serial_load_pre <= 1'b0;
                    if (serial_clock == 1'b0) begin
                        if (xfer_count == IO_CTRL_BITS - 1) begin
                            xfer_count <= 4'd0;
                            if (pad_count_2 == (19 + 19)) begin
                                xfer_state <= 2'b11;
                            end else begin
                                xfer_state <= 2'b01;
                            end
                        end else begin
                            xfer_count <= xfer_count + 1;
                        end
                    end else begin
                        serial_data_staging_1 <=
				{serial_data_staging_1[IO_CTRL_BITS-2:0], 1'b0};
                        serial_data_staging_2 <=
				{serial_data_staging_2[IO_CTRL_BITS-2:0], 1'b0};
                    end
		end
		2'b11: begin
                    xfer_count <= xfer_count + 1;

                    /* Load sequence:  Pulse clock for final data shift in;
                     * Pulse the load strobe.
                     * Return to idle mode.
                     */
                    if (xfer_count == 4'd0) begin
                        serial_clock_pre <= 1'b0;
                        serial_load_pre <= 1'b0;
                    end else if (xfer_count == 4'd1) begin
                        serial_clock_pre <= 1'b0;
                        serial_load_pre <= 1'b1;
                    end else if (xfer_count == 4'd2) begin
	    	    	serial_busy <= 1'b0;
                        serial_clock_pre <= 1'b0;
                        serial_load_pre <= 1'b0;
                        xfer_state <= 2'b00;
		    end
                end
            endcase
	end
    end

    // SPI Identification

    assign mfgr_id = 12'h456;		// Hard-coded
    assign prod_id = 8'h11;		// Hard-coded
    assign mask_rev = mask_rev_in;	// Copy in to out.

    // SPI Data transfer protocol.  The wishbone back door may only be
    // used if the front door is closed (CSB is high or the CSB pin is
    // not an input).  The time to apply values for the back door access
    // is limited to the clock cycle around the read or write from the
    // wbbd state machine (see below).

    assign caddr = (wbbd_busy) ? wbbd_addr : iaddr;
    assign csclk = (wbbd_busy) ? wbbd_sck : ((spi_is_active) ? mgmt_gpio_in[4] : 1'b0);
    assign cdata = (wbbd_busy) ? wbbd_data : idata;
    assign cwstb = (wbbd_busy) ? wbbd_write : wrstb;

    assign odata = fdata(caddr);

    // Register mapping and I/O to SPI interface module

    integer j;

    always @(posedge csclk or negedge porb) begin
	if (porb == 1'b0) begin
            // Set trim for PLL at (almost) slowest rate (~90MHz).  However,
            // pll_trim[12] must be set to zero for proper startup.
            pll_trim <= 26'b11111111111110111111111111;
            pll_sel <= 3'b010;		// Default output divider divide-by-2
            pll90_sel <= 3'b010;	// Default secondary output divider divide-by-2
            pll_div <= 5'b00100;	// Default feedback divider divide-by-8
            pll_dco_ena <= 1'b1;	// Default free-running PLL
            pll_ena <= 1'b0;		// Default PLL turned off
            pll_bypass <= 1'b1;		// Default bypass mode (don't use PLL)
            irq_spi <= 1'b0;
            reset_reg <= 1'b0;

	    // System monitoring signals
	    clk1_output_dest <= 1'b0;
	    clk2_output_dest <= 1'b0;
	    trap_output_dest <= 1'b0;
	    irq_1_inputsrc <= 1'b0;
	    irq_2_inputsrc <= 1'b0;

	    // GPIO Configuration, Data, and Control
	    // To-do:  Get user project pad defaults from external inputs
	    // to be configured by user or at project generation time.
	    // Pads 1 to 4 are the SPI and considered critical startup
	    // infrastructure, and should not be altered from the defaults
	    // below.  NOTE:  These are not startup values, but they should
	    // match the startup values applied to the GPIO, or else the
	    // GPIO should be always triggered to load at startup.

	    for (j = 0; j < (19 + 19); j=j+1) begin
		if ((j < 2) || (j >= (19 + 19) - 2)) begin
		    gpio_configure[j] <= 'h1803;
                end else begin
		    if (j == 3) begin
			// j == 3 corresponds to CSB, which is a weak pull-up
	                gpio_configure[j] <= 'h0801;
		    end else begin
	                gpio_configure[j] <= 'h0403;
		    end
		end
	    end

	    mgmt_gpio_data <= 'd0;
	    mgmt_gpio_data_buf <= 'd0;
	    serial_bb_enable <= 1'b0;
	    serial_bb_load <= 1'b0;
	    serial_bb_data_1 <= 1'b0;
	    serial_bb_data_2 <= 1'b0;
	    serial_bb_clock <= 1'b0;
	    serial_bb_resetn <= 1'b0;
	    serial_xfer <= 1'b0;
	    hkspi_disable <= 1'b0;
	    pwr_ctrl_out <= 'd0;







        end else begin
	    if (cwstb == 1'b1) begin
                case (caddr)
	    	    /* Register 8'h00 is reserved for future use */
	    	    /* Registers 8'h01 to 8'h07 are read-only and cannot be written */
            	    8'h08: begin
                	pll_ena <= cdata[0];
                	pll_dco_ena <= cdata[1];
            	    end
            	    8'h09: begin
                	pll_bypass <= cdata[0];
            	    end
            	    8'h0a: begin
                	irq_spi <= cdata[0];
            	    end
            	    8'h0b: begin
                	reset_reg <= cdata[0];
            	    end

		    /* Register 0c (trap state) is read-only */

            	    8'h0d: begin
                	pll_trim[7:0] <= cdata;
            	    end
            	    8'h0e: begin
                	pll_trim[15:8] <= cdata;
            	    end
            	    8'h0f: begin
                	pll_trim[23:16] <= cdata;
            	    end
            	    8'h10: begin
                	pll_trim[25:24] <= cdata[1:0];
            	    end
            	    8'h11: begin
                	pll90_sel <= cdata[5:3];
                	pll_sel <= cdata[2:0];
            	    end
            	    8'h12: begin
                	pll_div <= cdata[4:0];
            	    end
	    	    8'h13: begin
			serial_bb_data_2 <= cdata[6];
			serial_bb_data_1 <= cdata[5];
			serial_bb_clock  <= cdata[4];
			serial_bb_load   <= cdata[3];
			serial_bb_resetn <= cdata[2];
			serial_bb_enable <= cdata[1];
			serial_xfer <= cdata[0];
	    	    end











		    
		    /* Registers 16 to 19 (SRAM data) are read-only */

		    /* Register 1a (power monitor) is read-only */

            	    8'h1b: begin
			clk1_output_dest <= cdata[2];
			clk2_output_dest <= cdata[1];
			trap_output_dest <= cdata[0];
	    	    end
            	    8'h1c: begin
			irq_2_inputsrc <= cdata[1];
			irq_1_inputsrc <= cdata[0];
	    	    end
            	    8'h1d: begin
			gpio_configure[0][12:8] <= cdata[4:0];
	    	    end
            	    8'h1e: begin
			gpio_configure[0][7:0] <= cdata;
	    	    end
            	    8'h1f: begin
			gpio_configure[1][12:8] <= cdata[4:0];
	    	    end
            	    8'h20: begin
			gpio_configure[1][7:0] <= cdata;
	    	    end
            	    8'h21: begin
			gpio_configure[2][12:8] <= cdata[4:0];
	    	    end
            	    8'h22: begin
			gpio_configure[2][7:0] <= cdata;
	    	    end
            	    8'h23: begin
			gpio_configure[3][12:8] <= cdata[4:0];
	    	    end
            	    8'h24: begin
			gpio_configure[3][7:0] <= cdata;
	    	    end
            	    8'h25: begin
			gpio_configure[4][12:8] <= cdata[4:0];
	    	    end
            	    8'h26: begin
			gpio_configure[4][7:0] <= cdata;
	    	    end
            	    8'h27: begin
			gpio_configure[5][12:8] <= cdata[4:0];
	    	    end
            	    8'h28: begin
			gpio_configure[5][7:0] <= cdata;
	    	    end
            	    8'h29: begin
			gpio_configure[6][12:8] <= cdata[4:0];
	    	    end
            	    8'h2a: begin
			gpio_configure[6][7:0] <= cdata;
	    	    end
            	    8'h2b: begin
			gpio_configure[7][12:8] <= cdata[4:0];
	    	    end
            	    8'h2c: begin
			gpio_configure[7][7:0] <= cdata;
	    	    end
            	    8'h2d: begin
			gpio_configure[8][12:8] <= cdata[4:0];
	    	    end
            	    8'h2e: begin
			gpio_configure[8][7:0] <= cdata;
	    	    end
            	    8'h2f: begin
			gpio_configure[9][12:8] <= cdata[4:0];
	    	    end
            	    8'h30: begin
			gpio_configure[9][7:0] <= cdata;
	    	    end
            	    8'h31: begin
			gpio_configure[10][12:8] <= cdata[4:0];
	    	    end
            	    8'h32: begin
			gpio_configure[10][7:0] <= cdata;
	    	    end
            	    8'h33: begin
			gpio_configure[11][12:8] <= cdata[4:0];
	    	    end
            	    8'h34: begin
			gpio_configure[11][7:0] <= cdata;
	    	    end
            	    8'h35: begin
			gpio_configure[12][12:8] <= cdata[4:0];
	    	    end
            	    8'h36: begin
			gpio_configure[12][7:0] <= cdata;
	    	    end
            	    8'h37: begin
			gpio_configure[13][12:8] <= cdata[4:0];
	    	    end
            	    8'h38: begin
			gpio_configure[13][7:0] <= cdata;
	    	    end
            	    8'h39: begin
			gpio_configure[14][12:8] <= cdata[4:0];
	    	    end
            	    8'h3a: begin
			gpio_configure[14][7:0] <= cdata;
	    	    end
            	    8'h3b: begin
			gpio_configure[15][12:8] <= cdata[4:0];
	    	    end
            	    8'h3c: begin
			gpio_configure[15][7:0] <= cdata;
	    	    end
            	    8'h3d: begin
			gpio_configure[16][12:8] <= cdata[4:0];
	    	    end
            	    8'h3e: begin
			gpio_configure[16][7:0] <= cdata;
	    	    end
            	    8'h3f: begin
			gpio_configure[17][12:8] <= cdata[4:0];
	    	    end
            	    8'h40: begin
			gpio_configure[17][7:0] <= cdata;
	    	    end
            	    8'h41: begin
			gpio_configure[18][12:8] <= cdata[4:0];
	    	    end
            	    8'h42: begin
			gpio_configure[18][7:0] <= cdata;
	    	    end
            	    8'h43: begin
			gpio_configure[19][12:8] <= cdata[4:0];
	    	    end
            	    8'h44: begin
			gpio_configure[19][7:0] <= cdata;
	    	    end
            	    8'h45: begin
			gpio_configure[20][12:8] <= cdata[4:0];
	    	    end
            	    8'h46: begin
			gpio_configure[20][7:0] <= cdata;
	    	    end
            	    8'h47: begin
			gpio_configure[21][12:8] <= cdata[4:0];
	    	    end
            	    8'h48: begin
			gpio_configure[21][7:0] <= cdata;
	    	    end
            	    8'h49: begin
			gpio_configure[22][12:8] <= cdata[4:0];
	    	    end
            	    8'h4a: begin
			gpio_configure[22][7:0] <= cdata;
	    	    end
            	    8'h4b: begin
			gpio_configure[23][12:8] <= cdata[4:0];
	    	    end
            	    8'h4c: begin
			gpio_configure[23][7:0] <= cdata;
	    	    end
            	    8'h4d: begin
			gpio_configure[24][12:8] <= cdata[4:0];
	    	    end
            	    8'h4e: begin
			gpio_configure[24][7:0] <= cdata;
	    	    end
            	    8'h4f: begin
			gpio_configure[25][12:8] <= cdata[4:0];
	    	    end
            	    8'h50: begin
			gpio_configure[25][7:0] <= cdata;
	    	    end
            	    8'h51: begin
			gpio_configure[26][12:8] <= cdata[4:0];
	    	    end
            	    8'h52: begin
			gpio_configure[26][7:0] <= cdata;
	    	    end
            	    8'h53: begin
			gpio_configure[27][12:8] <= cdata[4:0];
	    	    end
            	    8'h54: begin
			gpio_configure[27][7:0] <= cdata;
	    	    end
            	    8'h55: begin
			gpio_configure[28][12:8] <= cdata[4:0];
	    	    end
            	    8'h56: begin
			gpio_configure[28][7:0] <= cdata;
	    	    end
            	    8'h57: begin
			gpio_configure[29][12:8] <= cdata[4:0];
	    	    end
            	    8'h58: begin
			gpio_configure[29][7:0] <= cdata;
	    	    end
            	    8'h59: begin
			gpio_configure[30][12:8] <= cdata[4:0];
	    	    end
            	    8'h5a: begin
			gpio_configure[30][7:0] <= cdata;
	    	    end
            	    8'h5b: begin
			gpio_configure[31][12:8] <= cdata[4:0];
	    	    end
            	    8'h5c: begin
			gpio_configure[31][7:0] <= cdata;
	    	    end
            	    8'h5d: begin
			gpio_configure[32][12:8] <= cdata[4:0];
	    	    end
            	    8'h5e: begin
			gpio_configure[32][7:0] <= cdata;
	    	    end
            	    8'h5f: begin
			gpio_configure[33][12:8] <= cdata[4:0];
	    	    end
            	    8'h60: begin
			gpio_configure[33][7:0] <= cdata;
	    	    end
            	    8'h61: begin
			gpio_configure[34][12:8] <= cdata[4:0];
	    	    end
            	    8'h62: begin
			gpio_configure[34][7:0] <= cdata;
	    	    end
            	    8'h63: begin
			gpio_configure[35][12:8] <= cdata[4:0];
	    	    end
            	    8'h64: begin
			gpio_configure[35][7:0] <= cdata;
	    	    end
            	    8'h65: begin
			gpio_configure[36][12:8] <= cdata[4:0];
	    	    end
            	    8'h66: begin
			gpio_configure[36][7:0] <= cdata;
	    	    end
            	    8'h67: begin
			gpio_configure[37][12:8] <= cdata[4:0];
	    	    end
            	    8'h68: begin
			gpio_configure[37][7:0] <= cdata;
	    	    end
	    	    8'h69: begin
			mgmt_gpio_data[37:32] <= cdata[5:0];
	    	    end
	    	    8'h6a: begin
			/* NOTE: mgmt_gpio_data updates only on the	*/
			/* upper byte write when writing through the	*/
			/* wishbone back-door.  This lets all bits	*/
			/* update at the same time.			*/
			if (spi_is_active) begin
			    mgmt_gpio_data[31:24] <= cdata;
			end else begin
			    mgmt_gpio_data[31:0] <= {cdata, mgmt_gpio_data_buf};
			end
	    	    end
	    	    8'h6b: begin
			if (spi_is_active) begin
			    mgmt_gpio_data[23:16] <= cdata;
			end else begin
			    mgmt_gpio_data_buf[23:16] <= cdata;
			end
	    	    end
	    	    8'h6c: begin
			if (spi_is_active) begin
			    mgmt_gpio_data[15:8] <= cdata;
			end else begin
			    mgmt_gpio_data_buf[15:8] <= cdata;
			end
	    	    end
	    	    8'h6d: begin
			if (spi_is_active) begin
			    mgmt_gpio_data[7:0] <= cdata;
			end else begin
			    mgmt_gpio_data_buf[7:0] <= cdata;
			end
	    	    end
	    	    8'h6e: begin
			pwr_ctrl_out <= cdata[3:0];
	    	    end
	    	    8'h6f: begin
			hkspi_disable <= cdata[0];
	    	    end
        	endcase	// (caddr)
    	    end else begin
	    	serial_xfer <= 1'b0;	// Serial transfer is self-resetting
		irq_spi <= 1'b0;	// IRQ is self-resetting
    	    end
    	end
    end
endmodule	// housekeeping

`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
// This routine synchronizes the 

module caravel_clocking(

    input VPWR,
    input VGND,

    input porb,		// Master (negative sense) reset from power-on-reset
    input resetb, 	// Master (negative sense) reset
    input ext_clk_sel,	// 0=use PLL clock, 1=use external (pad) clock
    input ext_clk,	// External pad (slow) clock
    input pll_clk,	// Internal PLL (fast) clock
    input pll_clk90,	// Internal PLL (fast) clock, 90 degree phase
    input [2:0] sel,	// Select clock divider value (0=thru, 1=divide-by-2, etc.)
    input [2:0] sel2,	// Select clock divider value for 90 degree phase divided clock
    input ext_reset,	// Positive sense reset from housekeeping SPI.
    output core_clk,	// Output core clock
    output user_clk,	// Output user (secondary) clock
    output resetb_sync	// Output propagated and buffered reset
);

    wire pll_clk_sel;
    wire pll_clk_divided;
    wire pll_clk90_divided;
    wire core_ext_clk;
    reg  use_pll_first;
    reg  use_pll_second;
    reg	 ext_clk_syncd_pre;
    reg	 ext_clk_syncd;

    wire resetb_async;

    assign pll_clk_sel = ~ext_clk_sel;

    assign resetb_async = porb & resetb & (!ext_reset);
    // Note that this implementation does not guard against switching to
    // the PLL clock if the PLL clock is not present.

    always @(posedge pll_clk or negedge resetb_async) begin
	if (resetb_async == 1'b0) begin
	    use_pll_first <= 1'b0;
	    use_pll_second <= 1'b0;
	    ext_clk_syncd <= 1'b0;
	end else begin
	    use_pll_first <= pll_clk_sel;
	    use_pll_second <= use_pll_first;
	    ext_clk_syncd_pre <= ext_clk;	// Sync ext_clk to pll_clk
	    ext_clk_syncd <= ext_clk_syncd_pre;	// Do this twice (resolve metastability)
	end
    end

    // Apply PLL clock divider

    clock_div #(
	.SIZE(3)
    ) divider (
	.in(pll_clk),
	.out(pll_clk_divided),
	.N(sel),
	.resetb(resetb_async)
    ); 

    // Secondary PLL clock divider for user space access

    clock_div #(
	.SIZE(3)
    ) divider2 (
	.in(pll_clk90),
	.out(pll_clk90_divided),
	.N(sel2),
	.resetb(resetb_async)
    ); 


    // Multiplex the clock output

    assign core_ext_clk = (use_pll_first) ? ext_clk_syncd : ext_clk;
    assign core_clk = (use_pll_second) ? pll_clk_divided : core_ext_clk;
    assign user_clk = (use_pll_second) ? pll_clk90_divided : core_ext_clk;

    // Reset assignment.  "reset" comes from POR, while "ext_reset"
    // comes from standalone SPI (and is normally zero unless
    // activated from the SPI).

    // Staged-delay reset
    reg [2:0] reset_delay;

    always @(negedge core_clk or negedge resetb_async) begin
        if (resetb_async == 1'b0) begin
        reset_delay <= 3'b111;
        end else begin
        reset_delay <= {1'b0, reset_delay[2:1]};
        end
    end

    assign resetb_sync = ~reset_delay[0];

endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
// Digital PLL (ring oscillator + controller)
// Technically this is a frequency locked loop, not a phase locked loop.






module digital_pll(

    VPWR,
    VGND,

    resetb, enable, osc, clockp, div, dco, ext_trim);


    input VPWR;
    input VGND;


    input	 resetb;	// Sense negative reset
    input	 enable;	// Enable PLL
    input	 osc;		// Input oscillator to match
    input [4:0]	 div;		// PLL feedback division ratio
    input 	 dco;		// Run in DCO mode
    input [25:0] ext_trim;	// External trim for DCO mode

    output [1:0] clockp;	// Two 90 degree clock phases

    wire [1:0]   clockp_buffer_in;	// Input wires to clockp buffers
    wire [25:0]  itrim;		// Internally generated trim bits
    wire [25:0]  otrim;		// Trim bits applied to the ring oscillator
    wire	 creset;	// Controller reset
    wire	 ireset;	// Internal reset (external reset OR disable)

    assign ireset = ~resetb | ~enable;

    // In DCO mode: Hold controller in reset and apply external trim value

    assign itrim = (dco == 1'b0) ? otrim : ext_trim;
    assign creset = (dco == 1'b0) ? ireset : 1'b1;

    (* keep *)
    ring_osc2x13 ringosc (
        .reset(ireset),
        .trim(itrim),
        .clockp(clockp_buffer_in)
    );

    digital_pll_controller pll_control (
        .reset(creset),
        .clock(clockp_buffer_in[0]),
        .osc(osc),
        .div(div),
        .trim(otrim)
    );

    (* keep *)
    sky130_fd_sc_hd__clkbuf_16 clockp_buffer_0 (

        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPWR),
        .VNB(VGND),

        .A(clockp_buffer_in[0]),
        .X(clockp[0])
    );

    (* keep *)
    sky130_fd_sc_hd__clkbuf_16 clockp_buffer_1 (

        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPWR),
        .VNB(VGND),

        .A(clockp_buffer_in[1]),
        .X(clockp[1])
    );

endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
// This module represents an unprogrammed mask revision
// block that is configured with via programming on the
// chip top level.  This value is passed to the block as
// a parameter

module user_id_programming #(
    parameter USER_PROJECT_ID = 32'h0
) (

    inout VPWR,
    inout VGND,

    output [31:0] mask_rev
);
    wire [31:0] user_proj_id_high;
    wire [31:0] user_proj_id_low;

    // For the mask revision input, use an array of digital constant logic cells

    sky130_fd_sc_hd__conb_1 mask_rev_value [31:0] (

            .VPWR(VPWR),
            .VPB(VPWR),
            .VNB(VGND),
            .VGND(VGND),

            .HI(user_proj_id_high),
            .LO(user_proj_id_low)
    );

    genvar i;
    generate
	for (i = 0; i < 32; i = i+1) begin
	    assign mask_rev[i] = (USER_PROJECT_ID & (32'h01 << i)) ?
			user_proj_id_high[i] : user_proj_id_low[i];
	end
    endgenerate

endmodule
`default_nettype wire
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module mprj_io_buffer (

      input VPWR,
      input VGND,

     input [(19-1):0]  mgmt_gpio_in,
     output [(19-1):0] mgmt_gpio_in_buf,
     input [2:0]   mgmt_gpio_oeb,
     output [2:0]  mgmt_gpio_oeb_buf,
     input [(19-1):0]  mgmt_gpio_out,
     output [(19-1):0] mgmt_gpio_out_buf
);


sky130_fd_sc_hd__clkbuf_8 BUF[(19*2+3)-1:0] (
    
            .VPWR(VPWR),
            .VGND(VGND),
            .VPB(VPWR),
            .VNB(VGND),
    
		.A({mgmt_gpio_in, mgmt_gpio_oeb, mgmt_gpio_out}), 
		.X({mgmt_gpio_in_buf, mgmt_gpio_oeb_buf, mgmt_gpio_out_buf})
); 

endmodulemodule buff_flash_clkrst (
	
		inout VPWR,
		inout VGND,
	
	input[11:0] in_n, 
	input[2:0] in_s, 
	output[11:0] out_s, 
	output[2:0] out_n);

	sky130_fd_sc_hd__clkbuf_8 BUF[14:0] (
		
			.VGND(VGND),
			.VNB(VGND),
			.VPB(VPWR),
			.VPWR(VPWR),
		
		.A({in_n, in_s}), 
		.X({out_s, out_n})); 

endmodule// SPDX-FileCopyrightText: 2022 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//	http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/*
 * gpio_signal_buffering ---
 *
 * This macro buffers long wires between housekeeping and the GPIO control
 * blocks at the top level of caravel.  The rule of thumb is to limit any
 * single wire length to approximately 1.3mm.  The physical (manhattan)
 * distances and required buffering are as follows:
 *
 * Breakpoints: 1.3, 2.6, 3.9, 5.2, 6.5, 7.8	(mm)
 * # buffers:     1,   2,   3,   4,   5,   6
 *
 * GPIO #    	wire length (mm)	# buffers
 *------------------------------------------------------
 * GPIO 0	0.4			0
 * GPIO 1	0.2			0
 * GPIO 2	0.0			0
 * GPIO 3	0.3			0
 * GPIO 4	0.5			0
 * GPIO 5	0.7			0
 * GPIO 6	1.0			0
 * GPIO 7	1.4			1	
 * GPIO 8	1.6			1
 * GPIO 9	1.8			1
 * GPIO 10	2.1			1
 * GPIO 11	2.3			1
 * GPIO 12	2.5			1
 * GPIO 13	2.7			2		
 * GPIO 14	3.6			2		
 * GPIO 15	4.5			3		
 * GPIO 16	4.7			3		
 * GPIO 17	5.1			3		
 * GPIO 18	5.4			4	   RHS
 *-------------------------------------------------------
 * GPIO 19	8.4			6	   LHS
 * GPIO 20	8.2			6
 * GPIO 21	7.9			6
 * GPIO 22	7.7			5
 * GPIO 23	7.4			5
 * GPIO 24	6.4			4
 * GPIO 25	6.1			4
 * GPIO 26	5.9			4
 * GPIO 27	5.7			4
 * GPIO 28	5.5			4
 * GPIO 29	5.3			4
 * GPIO 30	5.1			3
 * GPIO 31	4.8			3
 * GPIO 32	4.2			3
 * GPIO 33	4.0			3
 * GPIO 34	3.8			2
 * GPIO 35	3.5			2
 * GPIO 36	3.3			2
 * GPIO 37	3.4			2
 *------------------------------------------------------
 *	       total number of buffers: 95 (x2 for input and output)
 *
 * OEB lines go to GPIO 0 and 1 (no buffers needed) and GPIO 35-37
 * (2 buffers needed), so OEB lines need 6 additional buffers.
 *
 * The assumption is that all GPIOs on the left-hand side of the chip are
 * routed by taking wires left from the housekeeping across the top of the
 * SoC to the left side, and then up to the destination.  Right-hand side
 * connections go directly up the right side from the housekeeping block.
 *
 * Note that signal names are related to the signal being passed through;
 * "in" and "out" refer to the direction of the signal relative to the
 * housekeeping block in the top level.  For this macro, unbuffered signals
 * "unbuf" are the inputs, and buffered signals "buf" are the outputs.
 */

module gpio_signal_buffering (

	vccd,
	vssd,

    mgmt_io_in_unbuf,
    mgmt_io_out_unbuf,
    mgmt_io_oeb_buf,
    mgmt_io_in_buf,
    mgmt_io_out_buf,
    mgmt_io_oeb_unbuf
);


	input  vccd;
	input  vssd;


    /* NOTE:  To match the indices of the same signals in the
     * top level, add 35 to all OEB lines and add 7 to all in and out lines
     */
    input  [30:0] mgmt_io_in_unbuf;
    input  [30:0] mgmt_io_out_unbuf;
    input  [2:0] mgmt_io_oeb_unbuf;
    output [2:0] mgmt_io_oeb_buf;
    output [30:0] mgmt_io_in_buf;
    output [30:0] mgmt_io_out_buf;

    /* Instantiate 95 + 95 + 6 = 196 buffers of size 8 */

    wire [195:0] buf_in;
    wire [195:0] buf_out;

    sky130_fd_sc_hd__buf_8 signal_buffers [195:0] (
	
	    .VPWR(vccd),
	    .VGND(vssd),
	    .VPB(vccd),
	    .VNB(vssd),
	
	.A(buf_in),
	.X(buf_out)
    );

    /* Now chain them all together */

    //----------------------------------------
    // mgmt_io_in, right-hand side
    //----------------------------------------

    assign buf_in[0] = mgmt_io_in_unbuf[0];
    assign mgmt_io_in_buf[0] = buf_out[0];

    assign buf_in[1] = mgmt_io_in_unbuf[1];
    assign mgmt_io_in_buf[1] = buf_out[1];

    assign buf_in[2] = mgmt_io_in_unbuf[2];
    assign mgmt_io_in_buf[2] = buf_out[2];

    assign buf_in[3] = mgmt_io_in_unbuf[3];
    assign mgmt_io_in_buf[3] = buf_out[3];

    assign buf_in[4] = mgmt_io_in_unbuf[4];
    assign mgmt_io_in_buf[4] = buf_out[4];

    assign buf_in[5] = mgmt_io_in_unbuf[5];
    assign mgmt_io_in_buf[5] = buf_out[5];

    assign buf_in[6] = mgmt_io_in_unbuf[6];
    assign buf_in[7] = buf_out[6];
    assign mgmt_io_in_buf[6] = buf_out[7];

    assign buf_in[8] = mgmt_io_in_unbuf[7];
    assign buf_in[9] = buf_out[8];
    assign mgmt_io_in_buf[7] = buf_out[9];

    assign buf_in[10] = mgmt_io_in_unbuf[8];
    assign buf_in[11] = buf_out[10];
    assign buf_in[12] = buf_out[11];
    assign mgmt_io_in_buf[8] = buf_out[12];

    assign buf_in[13] = mgmt_io_in_unbuf[9];
    assign buf_in[14] = buf_out[13];
    assign buf_in[15] = buf_out[14];
    assign mgmt_io_in_buf[9] = buf_out[15];

    assign buf_in[16] = mgmt_io_in_unbuf[10];
    assign buf_in[17] = buf_out[16];
    assign buf_in[18] = buf_out[17];
    assign mgmt_io_in_buf[10] = buf_out[18];

    assign buf_in[19] = mgmt_io_in_unbuf[11];
    assign buf_in[20] = buf_out[19];
    assign buf_in[21] = buf_out[20];
    assign buf_in[22] = buf_out[21];
    assign mgmt_io_in_buf[11] = buf_out[22];

    //----------------------------------------
    // mgmt_io_in, left-hand side
    //----------------------------------------

    assign buf_in[23] = mgmt_io_in_unbuf[12];
    assign buf_in[24] = buf_out[23];
    assign buf_in[25] = buf_out[24];
    assign buf_in[26] = buf_out[25];
    assign buf_in[27] = buf_out[26];
    assign buf_in[28] = buf_out[27];
    assign mgmt_io_in_buf[12] = buf_out[28];

    assign buf_in[29] = mgmt_io_in_unbuf[13];
    assign buf_in[30] = buf_out[29];
    assign buf_in[31] = buf_out[30];
    assign buf_in[32] = buf_out[31];
    assign buf_in[33] = buf_out[32];
    assign buf_in[34] = buf_out[33];
    assign mgmt_io_in_buf[13] = buf_out[34];

    assign buf_in[35] = mgmt_io_in_unbuf[14];
    assign buf_in[36] = buf_out[35];
    assign buf_in[37] = buf_out[36];
    assign buf_in[38] = buf_out[37];
    assign buf_in[39] = buf_out[38];
    assign buf_in[40] = buf_out[39];
    assign mgmt_io_in_buf[14] = buf_out[40];

    assign buf_in[41] = mgmt_io_in_unbuf[15];
    assign buf_in[42] = buf_out[41];
    assign buf_in[43] = buf_out[42];
    assign buf_in[44] = buf_out[43];
    assign buf_in[45] = buf_out[44];
    assign mgmt_io_in_buf[15] = buf_out[45];

    assign buf_in[46] = mgmt_io_in_unbuf[16];
    assign buf_in[47] = buf_out[46];
    assign buf_in[48] = buf_out[47];
    assign buf_in[49] = buf_out[48];
    assign buf_in[50] = buf_out[49];
    assign mgmt_io_in_buf[16] = buf_out[50];

    assign buf_in[51] = mgmt_io_in_unbuf[17];
    assign buf_in[52] = buf_out[51];
    assign buf_in[53] = buf_out[52];
    assign buf_in[54] = buf_out[53];
    assign mgmt_io_in_buf[17] = buf_out[54];

    assign buf_in[55] = mgmt_io_in_unbuf[18];
    assign buf_in[56] = buf_out[55];
    assign buf_in[57] = buf_out[56];
    assign buf_in[58] = buf_out[57];
    assign mgmt_io_in_buf[18] = buf_out[58];

    assign buf_in[59] = mgmt_io_in_unbuf[19];
    assign buf_in[60] = buf_out[59];
    assign buf_in[61] = buf_out[60];
    assign buf_in[62] = buf_out[61];
    assign mgmt_io_in_buf[19] = buf_out[62];

    assign buf_in[63] = mgmt_io_in_unbuf[20];
    assign buf_in[64] = buf_out[63];
    assign buf_in[65] = buf_out[64];
    assign buf_in[66] = buf_out[65];
    assign mgmt_io_in_buf[20] = buf_out[66];

    assign buf_in[67] = mgmt_io_in_unbuf[21];
    assign buf_in[68] = buf_out[67];
    assign buf_in[69] = buf_out[68];
    assign buf_in[70] = buf_out[69];
    assign mgmt_io_in_buf[21] = buf_out[70];

    assign buf_in[71] = mgmt_io_in_unbuf[22];
    assign buf_in[72] = buf_out[71];
    assign buf_in[73] = buf_out[72];
    assign buf_in[74] = buf_out[73];
    assign mgmt_io_in_buf[22] = buf_out[74];

    assign buf_in[75] = mgmt_io_in_unbuf[23];
    assign buf_in[76] = buf_out[75];
    assign buf_in[77] = buf_out[76];
    assign mgmt_io_in_buf[23] = buf_out[77];

    assign buf_in[78] = mgmt_io_in_unbuf[24];
    assign buf_in[79] = buf_out[78];
    assign buf_in[80] = buf_out[79];
    assign mgmt_io_in_buf[24] = buf_out[80];

    assign buf_in[81] = mgmt_io_in_unbuf[25];
    assign buf_in[82] = buf_out[81];
    assign buf_in[83] = buf_out[82];
    assign mgmt_io_in_buf[25] = buf_out[83];

    assign buf_in[84] = mgmt_io_in_unbuf[26];
    assign buf_in[85] = buf_out[84];
    assign buf_in[86] = buf_out[85];
    assign mgmt_io_in_buf[26] = buf_out[86];

    assign buf_in[87] = mgmt_io_in_unbuf[27];
    assign buf_in[88] = buf_out[87];
    assign mgmt_io_in_buf[27] = buf_out[88];

    assign buf_in[89] = mgmt_io_in_unbuf[28];
    assign buf_in[90] = buf_out[89];
    assign mgmt_io_in_buf[28] = buf_out[90];

    assign buf_in[91] = mgmt_io_in_unbuf[29];
    assign buf_in[92] = buf_out[91];
    assign mgmt_io_in_buf[29] = buf_out[92];

    assign buf_in[93] = mgmt_io_in_unbuf[30];
    assign buf_in[94] = buf_out[93];
    assign mgmt_io_in_buf[30] = buf_out[94];

    //----------------------------------------
    // mgmt_io_out, right-hand side
    //----------------------------------------

    assign buf_in[95] = mgmt_io_out_unbuf[0];
    assign mgmt_io_out_buf[0] = buf_out[95];

    assign buf_in[96] = mgmt_io_out_unbuf[1];
    assign mgmt_io_out_buf[1] = buf_out[96];

    assign buf_in[97] = mgmt_io_out_unbuf[2];
    assign mgmt_io_out_buf[2] = buf_out[97];

    assign buf_in[98] = mgmt_io_out_unbuf[3];
    assign mgmt_io_out_buf[3] = buf_out[98];

    assign buf_in[99] = mgmt_io_out_unbuf[4];
    assign mgmt_io_out_buf[4] = buf_out[99];

    assign buf_in[100] = mgmt_io_out_unbuf[5];
    assign mgmt_io_out_buf[5] = buf_out[100];

    assign buf_in[101] = mgmt_io_out_unbuf[6];
    assign buf_in[102] = buf_out[101];
    assign mgmt_io_out_buf[6] = buf_out[102];

    assign buf_in[103] = mgmt_io_out_unbuf[7];
    assign buf_in[104] = buf_out[103];
    assign mgmt_io_out_buf[7] = buf_out[104];

    assign buf_in[105] = mgmt_io_out_unbuf[8];
    assign buf_in[106] = buf_out[105];
    assign buf_in[107] = buf_out[106];
    assign mgmt_io_out_buf[8] = buf_out[107];

    assign buf_in[108] = mgmt_io_out_unbuf[9];
    assign buf_in[109] = buf_out[108];
    assign buf_in[110] = buf_out[109];
    assign mgmt_io_out_buf[9] = buf_out[110];

    assign buf_in[111] = mgmt_io_out_unbuf[10];
    assign buf_in[112] = buf_out[111];
    assign buf_in[113] = buf_out[112];
    assign mgmt_io_out_buf[10] = buf_out[113];

    assign buf_in[114] = mgmt_io_out_unbuf[11];
    assign buf_in[115] = buf_out[114];
    assign buf_in[116] = buf_out[115];
    assign buf_in[117] = buf_out[116];
    assign mgmt_io_out_buf[11] = buf_out[117];

    //----------------------------------------
    // mgmt_io_out, left-hand side
    //----------------------------------------

    assign buf_in[118] = mgmt_io_out_unbuf[12];
    assign buf_in[119] = buf_out[118];
    assign buf_in[120] = buf_out[119];
    assign buf_in[121] = buf_out[120];
    assign buf_in[122] = buf_out[121];
    assign buf_in[123] = buf_out[122];
    assign mgmt_io_out_buf[12] = buf_out[123];

    assign buf_in[124] = mgmt_io_out_unbuf[13];
    assign buf_in[125] = buf_out[124];
    assign buf_in[126] = buf_out[125];
    assign buf_in[127] = buf_out[126];
    assign buf_in[128] = buf_out[127];
    assign buf_in[129] = buf_out[128];
    assign mgmt_io_out_buf[13] = buf_out[129];

    assign buf_in[130] = mgmt_io_out_unbuf[14];
    assign buf_in[131] = buf_out[130];
    assign buf_in[132] = buf_out[131];
    assign buf_in[133] = buf_out[132];
    assign buf_in[134] = buf_out[133];
    assign buf_in[135] = buf_out[134];
    assign mgmt_io_out_buf[14] = buf_out[135];

    assign buf_in[136] = mgmt_io_out_unbuf[15];
    assign buf_in[137] = buf_out[136];
    assign buf_in[138] = buf_out[137];
    assign buf_in[139] = buf_out[138];
    assign buf_in[140] = buf_out[139];
    assign mgmt_io_out_buf[15] = buf_out[140];

    assign buf_in[141] = mgmt_io_out_unbuf[16];
    assign buf_in[142] = buf_out[141];
    assign buf_in[143] = buf_out[142];
    assign buf_in[144] = buf_out[143];
    assign buf_in[145] = buf_out[144];
    assign mgmt_io_out_buf[16] = buf_out[145];

    assign buf_in[146] = mgmt_io_out_unbuf[17];
    assign buf_in[147] = buf_out[146];
    assign buf_in[148] = buf_out[147];
    assign buf_in[149] = buf_out[148];
    assign mgmt_io_out_buf[17] = buf_out[149];

    assign buf_in[150] = mgmt_io_out_unbuf[18];
    assign buf_in[151] = buf_out[150];
    assign buf_in[152] = buf_out[151];
    assign buf_in[153] = buf_out[152];
    assign mgmt_io_out_buf[18] = buf_out[153];

    assign buf_in[154] = mgmt_io_out_unbuf[19];
    assign buf_in[155] = buf_out[154];
    assign buf_in[156] = buf_out[155];
    assign buf_in[157] = buf_out[156];
    assign mgmt_io_out_buf[19] = buf_out[157];

    assign buf_in[158] = mgmt_io_out_unbuf[20];
    assign buf_in[159] = buf_out[158];
    assign buf_in[160] = buf_out[159];
    assign buf_in[161] = buf_out[160];
    assign mgmt_io_out_buf[20] = buf_out[161];

    assign buf_in[162] = mgmt_io_out_unbuf[21];
    assign buf_in[163] = buf_out[162];
    assign buf_in[164] = buf_out[163];
    assign buf_in[165] = buf_out[164];
    assign mgmt_io_out_buf[21] = buf_out[165];

    assign buf_in[166] = mgmt_io_out_unbuf[22];
    assign buf_in[167] = buf_out[166];
    assign buf_in[168] = buf_out[167];
    assign buf_in[169] = buf_out[168];
    assign mgmt_io_out_buf[22] = buf_out[169];

    assign buf_in[170] = mgmt_io_out_unbuf[23];
    assign buf_in[171] = buf_out[170];
    assign buf_in[172] = buf_out[171];
    assign mgmt_io_out_buf[23] = buf_out[172];

    assign buf_in[173] = mgmt_io_out_unbuf[24];
    assign buf_in[174] = buf_out[173];
    assign buf_in[175] = buf_out[174];
    assign mgmt_io_out_buf[24] = buf_out[175];

    assign buf_in[176] = mgmt_io_out_unbuf[25];
    assign buf_in[177] = buf_out[176];
    assign buf_in[178] = buf_out[177];
    assign mgmt_io_out_buf[25] = buf_out[178];

    assign buf_in[179] = mgmt_io_out_unbuf[26];
    assign buf_in[180] = buf_out[179];
    assign buf_in[181] = buf_out[180];
    assign mgmt_io_out_buf[26] = buf_out[181];

    assign buf_in[182] = mgmt_io_out_unbuf[27];
    assign buf_in[183] = buf_out[182];
    assign mgmt_io_out_buf[27] = buf_out[183];

    assign buf_in[184] = mgmt_io_out_unbuf[28];
    assign buf_in[185] = buf_out[184];
    assign mgmt_io_out_buf[28] = buf_out[185];

    assign buf_in[186] = mgmt_io_out_unbuf[29];
    assign buf_in[187] = buf_out[186];
    assign mgmt_io_out_buf[29] = buf_out[187];

    assign buf_in[188] = mgmt_io_out_unbuf[30];
    assign buf_in[189] = buf_out[188];
    assign mgmt_io_out_buf[30] = buf_out[189];

    //----------------------------------------
    // mgmt_io_oeb, left-hand side (only)
    //----------------------------------------

    assign buf_in[190] = mgmt_io_oeb_unbuf[0];
    assign buf_in[191] = buf_out[190];
    assign mgmt_io_oeb_buf[0] = buf_out[191];

    assign buf_in[192] = mgmt_io_oeb_unbuf[1];
    assign buf_in[193] = buf_out[192];
    assign mgmt_io_oeb_buf[1] = buf_out[193];

    assign buf_in[194] = mgmt_io_oeb_unbuf[2];
    assign buf_in[195] = buf_out[194];
    assign mgmt_io_oeb_buf[2] = buf_out[195];

  sky130_ef_sc_hd__decap_12 sigbuf_decaps [100:0] (
	
	    .VPWR(vccd),
	    .VGND(vssd),
	    .VPB(vccd),
	    .VNB(vssd)
	
  );

endmodule
 
 `default_nettype wire
 
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/*--------------------------------------------------------------*/
/* caravel, a project harness for the Google/SkyWater sky130	*/
/* fabrication process and open source PDK			*/
/*                                                          	*/
/* Copyright 2020 efabless, Inc.                            	*/
/* Written by Tim Edwards, December 2019                    	*/
/* and Mohamed Shalan, August 2020			    	*/
/* This file is open source hardware released under the     	*/
/* Apache 2.0 license.  See file LICENSE.                   	*/
/*								*/
/* Updated 10/15/2021:  Revised using the housekeeping module	*/
/* from housekeeping.v (refactoring a number of functions from	*/
/* the management SoC).						*/
/*                                                          	*/
/*--------------------------------------------------------------*/

module caravel_core (
    // All top-level I/O are package-facing pins

    inout vddio,  // Common 3.3V padframe/ESD power
    inout vssio,  // Common padframe/ESD ground
    inout vdda,   // Management 3.3V power
    inout vssa,   // Common analog ground
    inout vccd,   // Management/Common 1.8V power
    inout vssd,   // Common digital ground
    inout vdda1,  // User area 1 3.3V power
    inout vdda2,  // User area 2 3.3V power
    inout vssa1,  // User area 1 analog ground
    inout vssa2,  // User area 2 analog ground
    inout vccd1,  // User area 1 1.8V power
    inout vccd2,  // User area 2 1.8V power
    inout vssd1,  // User area 1 digital ground
    inout vssd2,  // User area 2 digital ground	


    // SoC Core Interface
    output porb_h,
    output por_l,
    input  rstb_h,
    input  clock_core,
    output gpio_out_core,
    input  gpio_in_core,
    output gpio_mode0_core,
    output gpio_mode1_core,
    output gpio_outenb_core,
    output gpio_inenb_core,

    // Flash SPI communication
    output flash_csb_frame,
    output flash_clk_frame,
    output flash_csb_oeb,
    output flash_clk_oeb,
    output flash_io0_oeb,
    output flash_io1_oeb,
    output flash_io0_ieb,
    output flash_io1_ieb,
    output flash_io0_do,
    output flash_io1_do,
    input  flash_io0_di,
    input  flash_io1_di,

    // User project IOs
    input  [  (19 + 19)-1:0] mprj_io_in,
    output [  (19 + 19)-1:0] mprj_io_out,
    output [  (19 + 19)-1:0] mprj_io_oeb,
    output [  (19 + 19)-1:0] mprj_io_inp_dis,
    output [  (19 + 19)-1:0] mprj_io_ib_mode_sel,
    output [  (19 + 19)-1:0] mprj_io_vtrip_sel,
    output [  (19 + 19)-1:0] mprj_io_slow_sel,
    output [  (19 + 19)-1:0] mprj_io_holdover,
    output [  (19 + 19)-1:0] mprj_io_analog_en,
    output [  (19 + 19)-1:0] mprj_io_analog_sel,
    output [  (19 + 19)-1:0] mprj_io_analog_pol,
    output [(19 + 19)*3-1:0] mprj_io_dm,

    // Loopbacks to constant value 1 in the 1.8V domain
    output [(19 + 19)-1:0] mprj_io_one,

    // User project direct access to gpio pad connections for analog
    // (all but the lowest-numbered 7 pads)
    inout [(19 + 19)-10:0] mprj_analog_io
);

    //------------------------------------------------------------
    // This value is uniquely defined for each user project.
    //------------------------------------------------------------
    parameter USER_PROJECT_ID = 32'h00000000;

    /*
     *--------------------------------------------------------------------
     *
     * These pins are overlaid on mprj_io space.  They have the function
     * below when the management processor is in reset, or in the default
     * configuration.  They are assigned to uses in the user space by the
     * configuration program running off of the SPI flash.  Note that even
     * when the user has taken control of these pins, they can be restored
     * to the original use by setting the resetb pin low.  The SPI pins and
     * UART pins can be connected directly to an FTDI chip as long as the
     * FTDI chip sets these lines to high impedence (input function) at
     * all times except when holding the chip in reset.
     *
     * JTAG       = mprj_io[0]		(inout)
     * SDO 	  = mprj_io[1]		(output)
     * SDI 	  = mprj_io[2]		(input)
     * CSB 	  = mprj_io[3]		(input)
     * SCK	  = mprj_io[4]		(input)
     * ser_rx     = mprj_io[5]		(input)
     * ser_tx     = mprj_io[6]		(output)
     * irq 	  = mprj_io[7]		(input)
     *
     * spi_sck    = mprj_io[32]		(output)
     * spi_csb    = mprj_io[33]		(output)
     * spi_sdi    = mprj_io[34]		(input)
     * spi_sdo    = mprj_io[35]		(output)
     * flash_io2  = mprj_io[36]		(inout) 
     * flash_io3  = mprj_io[37]		(inout) 
     *
     * These pins are reserved for any project that wants to incorporate
     * its own processor and flash controller.  While a user project can
     * technically use any available I/O pins for the purpose, these
     * four pins connect to a pass-through mode from the SPI slave (pins
     * 1-4 above) so that any SPI flash connected to these specific pins
     * can be accessed through the SPI slave even when the processor is in
     * reset.
     *
     * user_flash_csb = mprj_io[8]
     * user_flash_sck = mprj_io[9]
     * user_flash_io0 = mprj_io[10]
     * user_flash_io1 = mprj_io[11]
     *
     *--------------------------------------------------------------------
     */


    // User Project Control (user-facing)
    wire [(19 + 19)-1:0] user_io_oeb;
    wire [(19 + 19)-1:0] user_io_in;
    wire [(19 + 19)-1:0] user_io_out;

    /* Padframe control signals */
    wire [19-1:0] gpio_serial_link_1;
    wire [19-1:0] gpio_serial_link_2;
    wire mprj_io_loader_resetn;
    wire mprj_io_loader_clock;
    wire mprj_io_loader_strobe;
    wire mprj_io_loader_data_1;		/* user1 side serial loader */
    wire mprj_io_loader_data_2;		/* user2 side serial loader */

    // User Project Control management I/O
    // There are two types of GPIO connections:
    // (1) Full Bidirectional: Management connects to in, out, and oeb
    //     Uses:  JTAG and SDO
    // (2) Selectable bidirectional:  Management connects to in and out,
    //	   which are tied together.  oeb is grounded (oeb from the
    //	   configuration is used)

    // SDI 	 = mprj_io[2]		(input)
    // CSB 	 = mprj_io[3]		(input)
    // SCK	 = mprj_io[4]		(input)
    // ser_rx    = mprj_io[5]		(input)
    // ser_tx    = mprj_io[6]		(output)
    // irq 	 = mprj_io[7]		(input)

    wire [(19 + 19)-1:0] mgmt_io_in;	/* two- and three-pin data in	*/
    wire [(19 + 19)-1:0] mgmt_io_out;	/* two- and three-pin data out	*/
    wire [(19 + 19)-1:0] mgmt_io_oeb;	/* output enable, used only by	*/
						/* the three-pin interfaces	*/
    wire [(2 + 2)-1:0] pwr_ctrl_nc;	/* no-connects */

    // Power-on-reset signal.  The reset pad generates the sense-inverted
    // reset at 3.3V.  The 1.8V signal and the inverted 1.8V signal are
    // derived.
    wire rstb_l;

    // Flash SPI communication (management SoC to housekeeping)
    wire flash_clk_core,     flash_csb_core;
    wire flash_io0_oeb_core, flash_io1_oeb_core;
    wire flash_io2_oeb_core, flash_io3_oeb_core;
    wire flash_io0_ieb_core, flash_io1_ieb_core;
    wire flash_io2_ieb_core, flash_io3_ieb_core;
    wire flash_io0_do_core,  flash_io1_do_core;
    wire flash_io2_do_core,  flash_io3_do_core;
    wire flash_io0_di_core,  flash_io1_di_core;
    wire flash_io2_di_core,  flash_io3_di_core;


    // SoC core
    wire caravel_clk;
    wire caravel_clk2;
    wire caravel_rstn;

    // Logic analyzer signals
    wire [127:0] la_data_in_user;  // From CPU to MPRJ
    wire [127:0] la_data_in_mprj;  // From MPRJ to CPU
    wire [127:0] la_data_out_mprj; // From CPU to MPRJ
    wire [127:0] la_data_out_user; // From MPRJ to CPU
    wire [127:0] la_oenb_user;     // From CPU to MPRJ
    wire [127:0] la_oenb_mprj;     // From CPU to MPRJ
    wire [127:0] la_iena_mprj;     // From CPU only

    wire [2:0]   user_irq;	  // From MRPJ to CPU
    wire [2:0]   user_irq_core;
    wire [2:0]   user_irq_ena;
    wire [2:0]	 irq_spi;	  // From SPI and external pins

    // Exported Wishbone Bus (processor facing)
    wire mprj_iena_wb;
    wire mprj_cyc_o_core;
    wire mprj_stb_o_core;
    wire mprj_we_o_core;
    wire [3:0] mprj_sel_o_core;
    wire [31:0] mprj_adr_o_core;
    wire [31:0] mprj_dat_o_core;
    wire mprj_ack_i_core;
    wire [31:0] mprj_dat_i_core;

    wire [31:0] hk_dat_i;
    wire hk_ack_i;
    wire hk_stb_o;
    wire hk_cyc_o;

    // Exported Wishbone Bus (user area facing)
    wire 	mprj_cyc_o_user;
    wire 	mprj_stb_o_user;
    wire 	mprj_we_o_user;
    wire [3:0]  mprj_sel_o_user;
    wire [31:0] mprj_adr_o_user;
    wire [31:0] mprj_dat_o_user;
    wire [31:0] mprj_dat_i_user;
    wire	mprj_ack_i_user;

    // Mask revision
    wire [31:0] mask_rev;

    wire 	mprj_clock;
    wire 	mprj_clock2;
    wire 	mprj_reset;

    // Power monitoring 
    wire	mprj_vcc_pwrgood;
    wire	mprj2_vcc_pwrgood;
    wire	mprj_vdd_pwrgood;
    wire	mprj2_vdd_pwrgood;









    // Management processor (wrapper).  Any management core
    // implementation must match this pinout.

    mgmt_core_wrapper soc (
	
	    .VPWR(vccd),
	    .VGND(vssd),
	

	// Clock and reset
	.core_clk(caravel_clk),
	.core_rstn(caravel_rstn),

	// GPIO (1 pin)
	.gpio_out_pad(gpio_out_core),
	.gpio_in_pad(gpio_in_core),
	.gpio_mode0_pad(gpio_mode0_core),
	.gpio_mode1_pad(gpio_mode1_core),
	.gpio_outenb_pad(gpio_outenb_core),
	.gpio_inenb_pad(gpio_inenb_core),

	// Primary SPI flash controller
	.flash_csb(flash_csb_core),
	.flash_clk(flash_clk_core),
	.flash_io0_oeb(flash_io0_oeb_core),
	.flash_io0_di(flash_io0_di_core),
	.flash_io0_do(flash_io0_do_core),
	.flash_io1_oeb(flash_io1_oeb_core),
	.flash_io1_di(flash_io1_di_core),
	.flash_io1_do(flash_io1_do_core),
	.flash_io2_oeb(flash_io2_oeb_core),
	.flash_io2_di(flash_io2_di_core),
	.flash_io2_do(flash_io2_do_core),
	.flash_io3_oeb(flash_io3_oeb_core),
	.flash_io3_di(flash_io3_di_core),
	.flash_io3_do(flash_io3_do_core),

	// Exported Wishbone Bus
	.mprj_wb_iena(mprj_iena_wb),
	.mprj_cyc_o(mprj_cyc_o_core),
	.mprj_stb_o(mprj_stb_o_core),
	.mprj_we_o(mprj_we_o_core),
	.mprj_sel_o(mprj_sel_o_core),
	.mprj_adr_o(mprj_adr_o_core),
	.mprj_dat_o(mprj_dat_o_core),
	.mprj_ack_i(mprj_ack_i_core),
	.mprj_dat_i(mprj_dat_i_core),

	.hk_stb_o(hk_stb_o),
	.hk_cyc_o(hk_cyc_o),
	.hk_dat_i(hk_dat_i),
	.hk_ack_i(hk_ack_i),

	// IRQ
	.irq({irq_spi, user_irq}),
	.user_irq_ena(user_irq_ena),

	// Module status (these may or may not be implemented)
	.qspi_enabled(qspi_enabled),
	.uart_enabled(uart_enabled),
	.spi_enabled(spi_enabled),
	.debug_mode(debug_mode),

	// Module I/O (these may or may not be implemented)
	// UART
	.ser_tx(ser_tx),
	.ser_rx(ser_rx),
	// SPI master
	.spi_sdi(spi_sdi),
	.spi_csb(spi_csb),
	.spi_sck(spi_sck),
	.spi_sdo(spi_sdo),
	.spi_sdoenb(spi_sdoenb),
	// Debug
	.debug_in(debug_in),
	.debug_out(debug_out),
	.debug_oeb(debug_oeb),
	// Logic analyzer
	.la_input(la_data_in_mprj),
	.la_output(la_data_out_mprj),
	.la_oenb(la_oenb_mprj),
	.la_iena(la_iena_mprj),









	// Trap status
	.trap(trap)
    );

    /* Clock and reset to user space are passed through a tristate	*/
    /* buffer like the above, but since they are intended to be		*/
    /* always active, connect the enable to the logic-1 output from	*/
    /* the vccd1 domain.						*/

    mgmt_protect mgmt_buffers (
	
 	    .vccd(vccd),
	    .vssd(vssd),
	    .vccd1(vccd1),
	    .vssd1(vssd1),
	    .vccd2(vccd2),
	    .vssd2(vssd2),
	    .vdda1(vdda1),
	    .vssa1(vssa1),
	    .vdda2(vdda2),
	    .vssa2(vssa2),
	
	.caravel_clk(caravel_clk),
	.caravel_clk2(caravel_clk2),
	.caravel_rstn(caravel_rstn),

	.mprj_iena_wb(mprj_iena_wb),
	.mprj_cyc_o_core(mprj_cyc_o_core),
	.mprj_stb_o_core(mprj_stb_o_core),
	.mprj_we_o_core(mprj_we_o_core),
	.mprj_sel_o_core(mprj_sel_o_core),
	.mprj_adr_o_core(mprj_adr_o_core),
	.mprj_dat_o_core(mprj_dat_o_core),
	.mprj_ack_i_core(mprj_ack_i_core),
	.mprj_dat_i_core(mprj_dat_i_core),

	.user_irq_core(user_irq_core),
	.user_irq_ena(user_irq_ena),
	.la_data_out_core(la_data_out_user),
	.la_data_out_mprj(la_data_out_mprj),
	.la_data_in_core(la_data_in_user),
	.la_data_in_mprj(la_data_in_mprj),
	.la_oenb_mprj(la_oenb_mprj),
	.la_oenb_core(la_oenb_user),
	.la_iena_mprj(la_iena_mprj),

	.user_clock(mprj_clock),
	.user_clock2(mprj_clock2),
	.user_reset(mprj_reset),

	.mprj_cyc_o_user(mprj_cyc_o_user),
	.mprj_stb_o_user(mprj_stb_o_user),
	.mprj_we_o_user(mprj_we_o_user),
	.mprj_sel_o_user(mprj_sel_o_user),
	.mprj_adr_o_user(mprj_adr_o_user),
	.mprj_dat_o_user(mprj_dat_o_user),
	.mprj_dat_i_user(mprj_dat_i_user),
	.mprj_ack_i_user(mprj_ack_i_user),
	.user_irq(user_irq),
	.user1_vcc_powergood(mprj_vcc_pwrgood),
	.user2_vcc_powergood(mprj2_vcc_pwrgood),
	.user1_vdd_powergood(mprj_vdd_pwrgood),
	.user2_vdd_powergood(mprj2_vdd_pwrgood)
    );

    /*--------------------------------------------------*/
    /* Wrapper module around the user project 		*/
    /*--------------------------------------------------*/

    user_project_wrapper mprj ( 
        
	    .vdda1(vdda1),		// User area 1 3.3V power
	    .vdda2(vdda2),		// User area 2 3.3V power
	    .vssa1(vssa1),		// User area 1 analog ground
	    .vssa2(vssa2),		// User area 2 analog ground
	    .vccd1(vccd1),		// User area 1 1.8V power
	    .vccd2(vccd2),		// User area 2 1.8V power
	    .vssd1(vssd1),		// User area 1 digital ground
	    .vssd2(vssd2),		// User area 2 digital ground
    	

    	.wb_clk_i(mprj_clock),
    	.wb_rst_i(mprj_reset),

	// Management SoC Wishbone bus (exported)
	.wbs_cyc_i(mprj_cyc_o_user),
	.wbs_stb_i(mprj_stb_o_user),
	.wbs_we_i(mprj_we_o_user),
	.wbs_sel_i(mprj_sel_o_user),
	.wbs_adr_i(mprj_adr_o_user),
	.wbs_dat_i(mprj_dat_o_user),
	.wbs_ack_o(mprj_ack_i_user),
	.wbs_dat_o(mprj_dat_i_user),

	// GPIO pad 3-pin interface (plus analog)
	.io_in (user_io_in),
    .io_out(user_io_out),
    .io_oeb(user_io_oeb),
	.analog_io(mprj_analog_io),

	// Logic analyzer
	.la_data_in(la_data_in_user),
	.la_data_out(la_data_out_user),
	.la_oenb(la_oenb_user),

	// Independent clock
	.user_clock2(mprj_clock2),

	// IRQ
	.user_irq(user_irq_core)
    );

    /*------------------------------------------*/
    /* End user project instantiation		*/
    /*------------------------------------------*/

    wire [19-1:0] gpio_serial_link_1_shifted;
    wire [19-1:0] gpio_serial_link_2_shifted;

  assign gpio_serial_link_1_shifted = {
    gpio_serial_link_1[19-2:0], mprj_io_loader_data_1
  };
  // Note that serial_link_2 is backwards compared to serial_link_1, so it
  // shifts in the other direction.
  assign gpio_serial_link_2_shifted = {
    mprj_io_loader_data_2, gpio_serial_link_2[19-1:1]
  };

    // Propagating clock and reset to mitigate timing and fanout issues
    wire [19-1:0] gpio_clock_1;
    wire [19-1:0] gpio_clock_2;
    wire [19-1:0] gpio_resetn_1;
    wire [19-1:0] gpio_resetn_2;
    wire [19-1:0] gpio_load_1;
    wire [19-1:0] gpio_load_2;
    wire [19-1:0] gpio_clock_1_shifted;
    wire [19-1:0] gpio_clock_2_shifted;
    wire [19-1:0] gpio_resetn_1_shifted;
    wire [19-1:0] gpio_resetn_2_shifted;
    wire [19-1:0] gpio_load_1_shifted;
    wire [19-1:0] gpio_load_2_shifted;

  assign gpio_clock_1_shifted  = {gpio_clock_1[19-2:0], mprj_io_loader_clock};
  assign gpio_clock_2_shifted  = {mprj_io_loader_clock, gpio_clock_2[19-1:1]};
  assign gpio_resetn_1_shifted = {gpio_resetn_1[19-2:0], mprj_io_loader_resetn};
  assign gpio_resetn_2_shifted = {mprj_io_loader_resetn, gpio_resetn_2[19-1:1]};
  assign gpio_load_1_shifted   = {gpio_load_1[19-2:0], mprj_io_loader_strobe};
  assign gpio_load_2_shifted   = {mprj_io_loader_strobe, gpio_load_2[19-1:1]};

    wire [2:0] spi_pll_sel;
    wire [2:0] spi_pll90_sel;
    wire [4:0] spi_pll_div;
    wire [25:0] spi_pll_trim;

    // Clocking control

    caravel_clocking clock_ctrl (
    
		.VPWR(vccd),
		.VGND(vssd),
    
        .porb(porb_l),
        .ext_clk_sel(ext_clk_sel),
        .ext_clk(clock_core),
        .pll_clk(pll_clk),
        .pll_clk90(pll_clk90),
        .resetb(rstb_l),
        .sel(spi_pll_sel),
        .sel2(spi_pll90_sel),
        .ext_reset(ext_reset),  // From housekeeping SPI
        .core_clk(caravel_clk),
        .user_clk(caravel_clk2),
        .resetb_sync(caravel_rstn)
    );

    // DCO/Digital Locked Loop

    digital_pll pll (
    
		.VPWR(vccd),
		.VGND(vssd),
    
        .resetb(rstb_l),
        .enable(spi_pll_ena),
        .osc(clock_core),
        .clockp({pll_clk, pll_clk90}),
        .div(spi_pll_div),
        .dco(spi_pll_dco_ena),
        .ext_trim(spi_pll_trim)
    );


  // mprj_gpio_buffer signals
  wire [(19 + 19)-1:0] mgmt_io_in_hk;	/* mgmt_io_in at housekeeping	*/
  wire [(19 + 19)-1:0] mgmt_io_out_hk;	/* mgmt_io_out at housekeeping	*/
  wire [(19 + 19)-1:0] mgmt_io_oeb_hk;	/* mgmt_io_oeb at housekeeping	*/

  wire [(19-1):0] mgmt_gpio_in;
  wire [(19-1):0] mgmt_gpio_out;
  wire [2:0] mgmt_gpio_oeb;
  wire [(19-1):0] mgmt_gpio_in_buf;
  wire [(19-1):0] mgmt_gpio_out_buf;
  wire [2:0] mgmt_gpio_oeb_buf;

    // Housekeeping interface

    housekeeping housekeeping (
    
		.VPWR(vccd),
		.VGND(vssd),
    

        .wb_clk_i(caravel_clk),
        .wb_rstn_i(caravel_rstn),

        .wb_adr_i(mprj_adr_o_core),
        .wb_dat_i(mprj_dat_o_core),
        .wb_sel_i(mprj_sel_o_core),
        .wb_we_i(mprj_we_o_core),
        .wb_cyc_i(hk_cyc_o),
        .wb_stb_i(hk_stb_o),
        .wb_ack_o(hk_ack_i),
        .wb_dat_o(hk_dat_i),

        .porb(porb_l),

        .pll_ena(spi_pll_ena),
        .pll_dco_ena(spi_pll_dco_ena),
        .pll_div(spi_pll_div),
        .pll_sel(spi_pll_sel),
        .pll90_sel(spi_pll90_sel),
        .pll_trim(spi_pll_trim),
        .pll_bypass(ext_clk_sel),

	.qspi_enabled(qspi_enabled),
	.uart_enabled(uart_enabled),
	.spi_enabled(spi_enabled),
	.debug_mode(debug_mode),

	.ser_tx(ser_tx),
	.ser_rx(ser_rx),

	.spi_sdi(spi_sdi),
	.spi_csb(spi_csb),
	.spi_sck(spi_sck),
	.spi_sdo(spi_sdo),
	.spi_sdoenb(spi_sdoenb),

	.debug_in(debug_in),
	.debug_out(debug_out),
	.debug_oeb(debug_oeb),

        .irq(irq_spi),
        .reset(ext_reset),

        .serial_clock(mprj_io_loader_clock),
        .serial_load(mprj_io_loader_strobe),
        .serial_resetn(mprj_io_loader_resetn),
        .serial_data_1(mprj_io_loader_data_1),
        .serial_data_2(mprj_io_loader_data_2),

	.mgmt_gpio_in(mgmt_io_in_hk),
	.mgmt_gpio_out(mgmt_io_out_hk),
	.mgmt_gpio_oeb(mgmt_io_oeb_hk),

	.pwr_ctrl_out(pwr_ctrl_nc),	/* Not used in this version */

        .trap(trap),

	.user_clock(caravel_clk2),

        .mask_rev_in(mask_rev),

	.spimemio_flash_csb(flash_csb_core),
	.spimemio_flash_clk(flash_clk_core),
	.spimemio_flash_io0_oeb(flash_io0_oeb_core),
	.spimemio_flash_io1_oeb(flash_io1_oeb_core),
	.spimemio_flash_io2_oeb(flash_io2_oeb_core),
	.spimemio_flash_io3_oeb(flash_io3_oeb_core),
	.spimemio_flash_io0_do(flash_io0_do_core),
	.spimemio_flash_io1_do(flash_io1_do_core),
	.spimemio_flash_io2_do(flash_io2_do_core),
	.spimemio_flash_io3_do(flash_io3_do_core),
	.spimemio_flash_io0_di(flash_io0_di_core),
	.spimemio_flash_io1_di(flash_io1_di_core),
	.spimemio_flash_io2_di(flash_io2_di_core),
	.spimemio_flash_io3_di(flash_io3_di_core),

	.pad_flash_csb(flash_csb_frame),
	.pad_flash_csb_oeb(flash_csb_oeb),
	.pad_flash_clk(flash_clk_frame),
	.pad_flash_clk_oeb(flash_clk_oeb),
	.pad_flash_io0_oeb(flash_io0_oeb),
	.pad_flash_io1_oeb(flash_io1_oeb),
	.pad_flash_io0_ieb(flash_io0_ieb),
	.pad_flash_io1_ieb(flash_io1_ieb),
	.pad_flash_io0_do(flash_io0_do),
	.pad_flash_io1_do(flash_io1_do),
	.pad_flash_io0_di(flash_io0_di),
	.pad_flash_io1_di(flash_io1_di),








	.usr1_vcc_pwrgood(mprj_vcc_pwrgood),
	.usr2_vcc_pwrgood(mprj2_vcc_pwrgood),
	.usr1_vdd_pwrgood(mprj_vdd_pwrgood),
	.usr2_vdd_pwrgood(mprj2_vdd_pwrgood)
    );

  mprj_io_buffer gpio_buf (

      .VPWR(vccd),
      .VGND(vssd),


      .mgmt_gpio_in(mgmt_gpio_in),
      .mgmt_gpio_in_buf(mgmt_gpio_in_buf),
      .mgmt_gpio_oeb(mgmt_gpio_oeb),
      .mgmt_gpio_oeb_buf(mgmt_gpio_oeb_buf),
      .mgmt_gpio_out(mgmt_gpio_out),
      .mgmt_gpio_out_buf(mgmt_gpio_out_buf)
  );

  assign mgmt_gpio_in  = mgmt_io_in[((19 + 19)-1):(19)];
  assign mgmt_gpio_out = mgmt_io_out_hk[((19 + 19)-1):(19)];
  assign mgmt_gpio_oeb = mgmt_io_oeb_hk[((19 + 19)-1):((19 + 19)-3)];
  
  assign mgmt_io_in_hk = {mgmt_gpio_in_buf, mgmt_io_in[(19-1):0]};
  assign mgmt_io_out   = {mgmt_gpio_out_buf, mgmt_io_out_hk[(19-1):0]};
  assign mgmt_io_oeb   = {mgmt_gpio_oeb_buf, mgmt_io_oeb_hk[((19 + 19)-4):0]};

    /* GPIO defaults (via programmed) */
    wire [(19 + 19)*13-1:0] gpio_defaults;

    /* Fixed defaults for the first 5 GPIO pins */

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h1803)
    ) gpio_defaults_block_0 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[12:0])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h1803)
    ) gpio_defaults_block_1 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[25:13])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_2 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[38:26])
    );

    // CSB pin is set as an internal pull-up
    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0801)
    ) gpio_defaults_block_3 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[51:39])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_4 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[64:52])
    );

    /* Via-programmable defaults for the rest of the GPIO pins */

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_5 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[77:65])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_6 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[90:78])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_7 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[103:91])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_8 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[116:104])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_9 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[129:117])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_10 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[142:130])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_11 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[155:143])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_12 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[168:156])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_13 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[181:169])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_14 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[194:182])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_15 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[207:195])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_16 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[220:208])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_17 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[233:221])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_18 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[246:234])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_19 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[259:247])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_20 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[272:260])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_21 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[285:273])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_22 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[298:286])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_23 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[311:299])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_24 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[324:312])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_25 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[337:325])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_26 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[350:338])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_27 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[363:351])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_28 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[376:364])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_29 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[389:377])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_30 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[402:390])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_31 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[415:403])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_32 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[428:416])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_33 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[441:429])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_34 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[454:442])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_35 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[467:455])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_36 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[480:468])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_37 (
    	
	    .VPWR(vccd),
	    .VGND(vssd),
        
	.gpio_defaults(gpio_defaults[493:481])
    );

    // Each control block sits next to an I/O pad in the user area.
    // It gets input through a serial chain from the previous control
    // block and passes it to the next control block.  Due to the nature
    // of the shift register, bits are presented in reverse, as the first
    // bit in ends up as the last bit of the last I/O pad control block.

    // There are two types of block;  the first two and the last two
    // are configured to be full bidirectional under control of the
    // management Soc (JTAG and SDO for the first two;  flash_io2 and
    // flash_io3 for the last two).  The rest are configured to be default
    // (input).  Note that the first two and last two are the ones closest
    // to the management SoC on either side, which minimizes the wire length
    // of the extra signals those pads need.

    /* First two GPIOs (JTAG and SDO) */

    gpio_control_block gpio_control_bidir_1 [1:0] (
    	
	    .vccd(vccd),
	    .vssd(vssd),
	    .vccd1(vccd1),
	    .vssd1(vssd1),
        

	.gpio_defaults(gpio_defaults[25:0]),

    	// Management Soc-facing signals

    	.resetn(gpio_resetn_1_shifted[1:0]),
    	.serial_clock(gpio_clock_1_shifted[1:0]),
    	.serial_load(gpio_load_1_shifted[1:0]),

    	.resetn_out(gpio_resetn_1[1:0]),
    	.serial_clock_out(gpio_clock_1[1:0]),
    	.serial_load_out(gpio_load_1[1:0]),

    	.mgmt_gpio_in(mgmt_io_in[1:0]),
	.mgmt_gpio_out(mgmt_io_out[1:0]),
	.mgmt_gpio_oeb(mgmt_io_oeb[1:0]),

        .one(mprj_io_one[1:0]),
        .zero(),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_1_shifted[1:0]),
    	.serial_data_out(gpio_serial_link_1[1:0]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[1:0]),
    	.user_gpio_oeb(user_io_oeb[1:0]),
    	.user_gpio_in(user_io_in[1:0]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[1:0]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[1:0]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[1:0]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[1:0]),
    	.pad_gpio_holdover(mprj_io_holdover[1:0]),
    	.pad_gpio_ana_en(mprj_io_analog_en[1:0]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[1:0]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[1:0]),
    	.pad_gpio_dm(mprj_io_dm[5:0]),
    	.pad_gpio_outenb(mprj_io_oeb[1:0]),
    	.pad_gpio_out(mprj_io_out[1:0]),
    	.pad_gpio_in(mprj_io_in[1:0])
    );

    /* Section 1 GPIOs (GPIO 2 to 7) that start up under management control */

    gpio_control_block gpio_control_in_1a [5:0] (
        
            .vccd(vccd),
	    .vssd(vssd),
	    .vccd1(vccd1),
	    .vssd1(vssd1),
        

	.gpio_defaults(gpio_defaults[103:26]),

    	// Management Soc-facing signals

    	.resetn(gpio_resetn_1_shifted[7:2]),
    	.serial_clock(gpio_clock_1_shifted[7:2]),
    	.serial_load(gpio_load_1_shifted[7:2]),

    	.resetn_out(gpio_resetn_1[7:2]),
    	.serial_clock_out(gpio_clock_1[7:2]),
    	.serial_load_out(gpio_load_1[7:2]),

	.mgmt_gpio_in(mgmt_io_in[7:2]),
	.mgmt_gpio_out(mgmt_io_out[7:2]),
	.mgmt_gpio_oeb(mprj_io_one[7:2]),

        .one(mprj_io_one[7:2]),
        .zero(),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_1_shifted[7:2]),
    	.serial_data_out(gpio_serial_link_1[7:2]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[7:2]),
    	.user_gpio_oeb(user_io_oeb[7:2]),
    	.user_gpio_in(user_io_in[7:2]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[7:2]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[7:2]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[7:2]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[7:2]),
    	.pad_gpio_holdover(mprj_io_holdover[7:2]),
    	.pad_gpio_ana_en(mprj_io_analog_en[7:2]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[7:2]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[7:2]),
    	.pad_gpio_dm(mprj_io_dm[23:6]),
    	.pad_gpio_outenb(mprj_io_oeb[7:2]),
    	.pad_gpio_out(mprj_io_out[7:2]),
    	.pad_gpio_in(mprj_io_in[7:2])
    );

    /* Section 1 GPIOs (GPIO 8 to 18) */

    gpio_control_block gpio_control_in_1 [19-9:0] (
        
            .vccd(vccd),
	    .vssd(vssd),
	    .vccd1(vccd1),
	    .vssd1(vssd1),
        

	.gpio_defaults(gpio_defaults[(19*13-1):104]),

    	// Management Soc-facing signals

    	.resetn(gpio_resetn_1_shifted[(19-1):8]),
    	.serial_clock(gpio_clock_1_shifted[(19-1):8]),
    	.serial_load(gpio_load_1_shifted[(19-1):8]),

    	.resetn_out(gpio_resetn_1[(19-1):8]),
    	.serial_clock_out(gpio_clock_1[(19-1):8]),
    	.serial_load_out(gpio_load_1[(19-1):8]),

	.mgmt_gpio_in(mgmt_io_in[(19-1):8]),
	.mgmt_gpio_out(mgmt_io_out[(19-1):8]),
	.mgmt_gpio_oeb(mprj_io_one[(19-1):8]),
  
        .one(mprj_io_one[(19-1):8]),
        .zero(),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_1_shifted[(19-1):8]),
    	.serial_data_out(gpio_serial_link_1[(19-1):8]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[(19-1):8]),
    	.user_gpio_oeb(user_io_oeb[(19-1):8]),
    	.user_gpio_in(user_io_in[(19-1):8]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[(19-1):8]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[(19-1):8]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[(19-1):8]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[(19-1):8]),
    	.pad_gpio_holdover(mprj_io_holdover[(19-1):8]),
    	.pad_gpio_ana_en(mprj_io_analog_en[(19-1):8]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[(19-1):8]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[(19-1):8]),
    	.pad_gpio_dm(mprj_io_dm[(19*3-1):24]),
    	.pad_gpio_outenb(mprj_io_oeb[(19-1):8]),
    	.pad_gpio_out(mprj_io_out[(19-1):8]),
    	.pad_gpio_in(mprj_io_in[(19-1):8])
    );

    /* Last three GPIOs (spi_sdo, flash_io2, and flash_io3) */

    gpio_control_block gpio_control_bidir_2 [2:0] (
    	
	    .vccd(vccd),
	    .vssd(vssd),
	    .vccd1(vccd1),
	    .vssd1(vssd1),
        

	.gpio_defaults(gpio_defaults[((19 + 19)*13-1):((19 + 19)*13-39)]),

    	// Management Soc-facing signals

    	.resetn(gpio_resetn_2_shifted[(19-1):(19-3)]),
    	.serial_clock(gpio_clock_2_shifted[(19-1):(19-3)]),
    	.serial_load(gpio_load_2_shifted[(19-1):(19-3)]),

    	.resetn_out(gpio_resetn_2[(19-1):(19-3)]),
    	.serial_clock_out(gpio_clock_2[(19-1):(19-3)]),
    	.serial_load_out(gpio_load_2[(19-1):(19-3)]),

    	.mgmt_gpio_in(mgmt_io_in[((19 + 19)-1):((19 + 19)-3)]),
	.mgmt_gpio_out(mgmt_io_out[((19 + 19)-1):((19 + 19)-3)]),
	.mgmt_gpio_oeb(mgmt_io_oeb[((19 + 19)-1):((19 + 19)-3)]),

        .one(mprj_io_one[((19 + 19)-1):((19 + 19)-3)]),
        .zero(),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_2_shifted[(19-1):(19-3)]),
    	.serial_data_out(gpio_serial_link_2[(19-1):(19-3)]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[((19 + 19)-1):((19 + 19)-3)]),
    	.user_gpio_oeb(user_io_oeb[((19 + 19)-1):((19 + 19)-3)]),
    	.user_gpio_in(user_io_in[((19 + 19)-1):((19 + 19)-3)]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_holdover(mprj_io_holdover[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_ana_en(mprj_io_analog_en[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_dm(mprj_io_dm[((19 + 19)*3-1):((19 + 19)*3-9)]),
    	.pad_gpio_outenb(mprj_io_oeb[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_out(mprj_io_out[((19 + 19)-1):((19 + 19)-3)]),
    	.pad_gpio_in(mprj_io_in[((19 + 19)-1):((19 + 19)-3)])
    );

    /* Section 2 GPIOs (GPIO 19 to 34) */

    gpio_control_block gpio_control_in_2 [19-4:0] (
    	
            .vccd(vccd),
	    .vssd(vssd),
	    .vccd1(vccd1),
	    .vssd1(vssd1),
        

	.gpio_defaults(gpio_defaults[((19 + 19)*13-40):(19*13)]),

    	// Management Soc-facing signals

    	.resetn(gpio_resetn_2_shifted[(19-4):0]),
    	.serial_clock(gpio_clock_2_shifted[(19-4):0]),
    	.serial_load(gpio_load_2_shifted[(19-4):0]),

    	.resetn_out(gpio_resetn_2[(19-4):0]),
    	.serial_clock_out(gpio_clock_2[(19-4):0]),
    	.serial_load_out(gpio_load_2[(19-4):0]),

	.mgmt_gpio_in(mgmt_io_in[((19 + 19)-4):(19)]),
	.mgmt_gpio_out(mgmt_io_out[((19 + 19)-4):(19)]),
	.mgmt_gpio_oeb(mprj_io_one[((19 + 19)-4):(19)]),


        .one(mprj_io_one[((19 + 19)-4):(19)]),
        .zero(),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_2_shifted[(19-4):0]),
    	.serial_data_out(gpio_serial_link_2[(19-4):0]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[((19 + 19)-4):(19)]),
    	.user_gpio_oeb(user_io_oeb[((19 + 19)-4):(19)]),
    	.user_gpio_in(user_io_in[((19 + 19)-4):(19)]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[((19 + 19)-4):(19)]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[((19 + 19)-4):(19)]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[((19 + 19)-4):(19)]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[((19 + 19)-4):(19)]),
    	.pad_gpio_holdover(mprj_io_holdover[((19 + 19)-4):(19)]),
    	.pad_gpio_ana_en(mprj_io_analog_en[((19 + 19)-4):(19)]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[((19 + 19)-4):(19)]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[((19 + 19)-4):(19)]),
    	.pad_gpio_dm(mprj_io_dm[((19 + 19)*3-10):(19*3)]),
    	.pad_gpio_outenb(mprj_io_oeb[((19 + 19)-4):(19)]),
    	.pad_gpio_out(mprj_io_out[((19 + 19)-4):(19)]),
    	.pad_gpio_in(mprj_io_in[((19 + 19)-4):(19)])
    );

    user_id_programming #(
	.USER_PROJECT_ID(USER_PROJECT_ID)
    ) user_id_value (
	
		.VPWR(vccd),
		.VGND(vssd),
	
	.mask_rev(mask_rev)
    );

    // Power-on-reset circuit
    simple_por por (
	
		.vdd3v3(vddio),
		.vdd1v8(vccd),
		.vss3v3(vssio),
		.vss1v8(vssd),
	
		.porb_h(porb_h),
		.porb_l(porb_l),
		.por_l(por_l)
    );

    // XRES (chip input pin reset) reset level converter
    xres_buf rstb_level (
	
		.VPWR(vddio),
		.LVPWR(vccd),
		.LVGND(vssd),
		.VGND(vssio),
	
		.A(rstb_h),
		.X(rstb_l)
    );

    /* Spare logic for metal mask fixes */
    // `define NUM_SPARE_BLOCKS (`MPRJ_IO_PADS+4)
    

    wire [(27*4)-1:0] spare_xz_nc;
    wire [(4*4)-1:0] spare_xi_nc;
    wire [(1*4)-1:0] spare_xib_nc;
    wire [(2*4)-1:0] spare_xna_nc;
    wire [(2*4)-1:0] spare_xno_nc;
    wire [(2*4)-1:0] spare_xmx_nc;
    wire [(2*4)-1:0] spare_xfq_nc;
    wire [(2*4)-1:0] spare_xfqn_nc;

    // Four spare logic blocks above the processor and one per GPIO
    // control block.
(* keep *) spare_logic_block spare_logic [4-1:0] (
	
		.vccd(vccd),
		.vssd(vssd),
	
		.spare_xz(spare_xz_nc),
		.spare_xi(spare_xi_nc),
		.spare_xib(spare_xib_nc),
		.spare_xna(spare_xna_nc),
		.spare_xno(spare_xno_nc),
		.spare_xmx(spare_xmx_nc),
		.spare_xfq(spare_xfq_nc),
		.spare_xfqn(spare_xfqn_nc)
    );
(* keep *) empty_macro empty_macro_0 ();
(* keep *) empty_macro empty_macro_1 ();
(* keep *) manual_power_connections manual_power_connections ();
endmodule
// `default_nettype wire 
 `default_nettype wire
 
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/*--------------------------------------------------------------*/
/* caravel, a project harness for the Google/SkyWater sky130	*/
/* fabrication process and open source PDK			*/
/*                                                          	*/
/* Copyright 2020 efabless, Inc.                            	*/
/* Written by Tim Edwards, December 2019                    	*/
/* and Mohamed Shalan, August 2020			    	*/
/* This file is open source hardware released under the     	*/
/* Apache 2.0 license.  See file LICENSE.                   	*/
/*								*/
/* Updated 10/15/2021:  Revised using the housekeeping module	*/
/* from housekeeping.v (refactoring a number of functions from	*/
/* the management SoC).						*/
/*                                                          	*/
/*--------------------------------------------------------------*/

module caravel (
    // All top-level I/O are package-facing pins
    inout                     vddio,    // Common 3.3V padframe/ESD power
    inout                     vddio_2,  // Common 3.3V padframe/ESD power
    inout                     vssio,    // Common padframe/ESD ground
    inout                     vssio_2,  // Common padframe/ESD ground
    inout                     vdda,     // Management 3.3V power
    inout                     vssa,     // Common analog ground
    inout                     vccd,     // Management/Common 1.8V power
    inout                     vssd,     // Common digital ground
    inout                     vdda1,    // User area 1 3.3V power
    inout                     vdda1_2,  // User area 1 3.3V power
    inout                     vdda2,    // User area 2 3.3V power
    inout                     vssa1,    // User area 1 analog ground
    inout                     vssa1_2,  // User area 1 analog ground
    inout                     vssa2,    // User area 2 analog ground
    inout                     vccd1,    // User area 1 1.8V power
    inout                     vccd2,    // User area 2 1.8V power
    inout                     vssd1,    // User area 1 digital ground
    inout                     vssd2,    // User area 2 digital ground	
    inout                     gpio,     // Used for external LDO control
    inout [(19 + 19)-1:0] mprj_io,
    input                     clock,    // CMOS core clock input, not a crystal
    input                     resetb,   // Reset input (Active Low)

    // Note that only two flash data pins are dedicated to the
    // management SoC wrapper.  The management SoC exports the
    // quad SPI mode status to make use of the top two mprj_io
    // pins for io2 and io3.
    output flash_csb,
    output flash_clk,
    inout  flash_io0,
    inout  flash_io1
);

  //------------------------------------------------------------
  // This value is uniquely defined for each user project.
  //------------------------------------------------------------
  parameter USER_PROJECT_ID = 32'h00000000;

  /*
     *--------------------------------------------------------------------
     * These pins are overlaid on mprj_io space. They have the function
     * below when the management processor is in reset, or in the default
     * configuration. They are assigned to uses in the user space by the
     * configuration program running off of the SPI flash.  Note that even
     * when the user has taken control of these pins, they can be restored
     * to the original use by setting the resetb pin low.  The SPI pins and
     * UART pins can be connected directly to an FTDI chip as long as the
     * FTDI chip sets these lines to high impedence (input function) at
     * all times except when holding the chip in reset.
     *
     * JTAG			= mprj_io[0]		(inout)
     * SDO			= mprj_io[1]		(output)
     * SDI			= mprj_io[2]		(input)
     * CSB			= mprj_io[3]		(input)
     * SCK			= mprj_io[4]		(input)
     * ser_rx		= mprj_io[5]		(input)
     * ser_tx		= mprj_io[6]		(output)
     * irq			= mprj_io[7]		(input)
     *
     * spi_sck		= mprj_io[32]		(output)
     * spi_csb		= mprj_io[33]		(output)
     * spi_sdi		= mprj_io[34]		(input)
     * spi_sdo		= mprj_io[35]		(output)
     * flash_io2	= mprj_io[36]		(inout) 
     * flash_io3	= mprj_io[37]		(inout) 
     *
     * These pins are reserved for any project that wants to incorporate
     * its own processor and flash controller.  While a user project can
     * technically use any available I/O pins for the purpose, these
     * four pins connect to a pass-through mode from the SPI slave (pins
     * 1-4 above) so that any SPI flash connected to these specific pins
     * can be accessed through the SPI slave even when the processor is in
     * reset.
     *
     * user_flash_csb = mprj_io[8]
     * user_flash_sck = mprj_io[9]
     * user_flash_io0 = mprj_io[10]
     * user_flash_io1 = mprj_io[11]
     *
     *--------------------------------------------------------------------
     */

  // One-bit GPIO dedicated to management SoC (outside of user control)
  wire gpio_out_core;
  wire gpio_in_core;
  wire gpio_mode0_core;
  wire gpio_mode1_core;
  wire gpio_outenb_core;
  wire gpio_inenb_core;

  // User Project Control (pad-facing)
  wire [(19 + 19)-1:0] mprj_io_inp_dis;
  wire [(19 + 19)-1:0] mprj_io_oeb;
  wire [(19 + 19)-1:0] mprj_io_ib_mode_sel;
  wire [(19 + 19)-1:0] mprj_io_vtrip_sel;
  wire [(19 + 19)-1:0] mprj_io_slow_sel;
  wire [(19 + 19)-1:0] mprj_io_holdover;
  wire [(19 + 19)-1:0] mprj_io_analog_en;
  wire [(19 + 19)-1:0] mprj_io_analog_sel;
  wire [(19 + 19)-1:0] mprj_io_analog_pol;
  wire [(19 + 19)*3-1:0] mprj_io_dm;
  wire [(19 + 19)-1:0] mprj_io_in;
  wire [(19 + 19)-1:0] mprj_io_out;
  wire [(19 + 19)-1:0] mprj_io_one;

  // User Project Control (user-facing)
  wire [(19 + 19)-10:0] user_analog_io;

  // User Project Control management I/O
  // There are two types of GPIO connections:
  // (1) Full Bidirectional: Management connects to in, out, and oeb
  //     Uses:  JTAG and SDO
  // (2) Selectable bidirectional:  Management connects to in and out,
  //	   which are tied together.  oeb is grounded (oeb from the
  //	   configuration is used)

  // SDI		= mprj_io[2]		(input)
  // CSB		= mprj_io[3]		(input)
  // SCK		= mprj_io[4]		(input)
  // ser_rx	= mprj_io[5]		(input)
  // ser_tx	= mprj_io[6]		(output)
  // irq		= mprj_io[7]		(input)

  wire clock_core;

  // Power-on-reset signal.  The reset pad generates the sense-inverted
  // reset at 3.3V.  The 1.8V signal and the inverted 1.8V signal are
  // derived.

  wire porb_h;
  wire porb_l;
  wire por_l;

  wire rstb_h;

  // Flash SPI communication (
  wire flash_clk_frame;
  wire flash_csb_frame;
  wire flash_clk_oeb, flash_csb_oeb;
  wire flash_clk_ieb, flash_csb_ieb;
  wire flash_io0_oeb, flash_io1_oeb;
  wire flash_io0_ieb, flash_io1_ieb;
  wire flash_io0_do, flash_io1_do;
  wire flash_io0_di, flash_io1_di;

  wire vddio_core;
  wire vssio_core;
  wire vdda_core;
  wire vssa_core;
  wire vccd_core;
  wire vssd_core;
  wire vdda1_core;
  wire vdda2_core;
  wire vssa1_core;
  wire vssa2_core;
  wire vccd1_core;
  wire vccd2_core;
  wire vssd1_core;
  wire vssd2_core;

  chip_io padframe (

      // Package Pins
      .vddio_pad(vddio),  // Common padframe/ESD supply
      .vddio_pad2(vddio_2),
      .vssio_pad(vssio),  // Common padframe/ESD ground
      .vssio_pad2(vssio_2),
      .vccd_pad(vccd),  // Common 1.8V supply
      .vssd_pad(vssd),  // Common digital ground
      .vdda_pad(vdda),  // Management analog 3.3V supply
      .vssa_pad(vssa),  // Management analog ground
      .vdda1_pad(vdda1),  // User area 1 3.3V supply
      .vdda1_pad2(vdda1_2),
      .vdda2_pad(vdda2),  // User area 2 3.3V supply
      .vssa1_pad(vssa1),  // User area 1 analog ground
      .vssa1_pad2(vssa1_2),
      .vssa2_pad(vssa2),  // User area 2 analog ground
      .vccd1_pad(vccd1),  // User area 1 1.8V supply
      .vccd2_pad(vccd2),  // User area 2 1.8V supply
      .vssd1_pad(vssd1),  // User area 1 digital ground
      .vssd2_pad(vssd2),  // User area 2 digital ground
      .vddio(vddio_core),
      .vssio(vssio_core),
      .vdda(vdda_core),
      .vssa(vssa_core),
      .vccd(vccd_core),
      .vssd(vssd_core),
      .vdda1(vdda1_core),
      .vdda2(vdda2_core),
      .vssa1(vssa1_core),
      .vssa2(vssa2_core),
      .vccd1(vccd1_core),
      .vccd2(vccd2_core),
      .vssd1(vssd1_core),
      .vssd2(vssd2_core),
      
      // Core Side Pins
      .gpio(gpio),
      .mprj_io(mprj_io),
      .clock(clock),
      .resetb(resetb),
      .flash_csb(flash_csb),
      .flash_clk(flash_clk),
      .flash_io0(flash_io0),
      .flash_io1(flash_io1),


      // SoC Core Interface
      .porb_h(porb_h),
      .por(por_l),
      .resetb_core_h(rstb_h),
      .clock_core(clock_core),
      .gpio_out_core(gpio_out_core),
      .gpio_in_core(gpio_in_core),
      .gpio_mode0_core(gpio_mode0_core),
      .gpio_mode1_core(gpio_mode1_core),
      .gpio_outenb_core(gpio_outenb_core),
      .gpio_inenb_core(gpio_inenb_core),
      .flash_csb_core(flash_csb_frame),
      .flash_clk_core(flash_clk_frame),
      .flash_csb_oeb_core(flash_csb_oeb),
      .flash_clk_oeb_core(flash_clk_oeb),
      .flash_io0_oeb_core(flash_io0_oeb),
      .flash_io1_oeb_core(flash_io1_oeb),
      .flash_io0_ieb_core(flash_io0_ieb),
      .flash_io1_ieb_core(flash_io1_ieb),
      .flash_io0_do_core(flash_io0_do),
      .flash_io1_do_core(flash_io1_do),
      .flash_io0_di_core(flash_io0_di),
      .flash_io1_di_core(flash_io1_di),
      .mprj_io_one(mprj_io_one),
      .mprj_io_in(mprj_io_in),
      .mprj_io_out(mprj_io_out),
      .mprj_io_oeb(mprj_io_oeb),
      .mprj_io_inp_dis(mprj_io_inp_dis),
      .mprj_io_ib_mode_sel(mprj_io_ib_mode_sel),
      .mprj_io_vtrip_sel(mprj_io_vtrip_sel),
      .mprj_io_slow_sel(mprj_io_slow_sel),
      .mprj_io_holdover(mprj_io_holdover),
      .mprj_io_analog_en(mprj_io_analog_en),
      .mprj_io_analog_sel(mprj_io_analog_sel),
      .mprj_io_analog_pol(mprj_io_analog_pol),
      .mprj_io_dm(mprj_io_dm),
      .mprj_analog_io(user_analog_io)
  );

  caravel_core chip_core (
      // All top-level I/O are package-facing pins

      .vddio(vddio_core),  // Common 3.3V padframe/ESD power
      .vssio(vssio_core),  // Common padframe/ESD ground
//    .vdda (vdda_core),   // Management 3.3V power
//    .vssa (vssa_core),   // Common analog ground
      .vccd (vccd_core),   // Management/Common 1.8V power
      .vssd (vssd_core),   // Common digital ground
      .vdda1(vdda1_core),  // User area 1 3.3V power
      .vdda2(vdda2_core),  // User area 2 3.3V power
      .vssa1(vssa1_core),  // User area 1 analog ground
      .vssa2(vssa2_core),  // User area 2 analog ground
      .vccd1(vccd1_core),  // User area 1 1.8V power
      .vccd2(vccd2_core),  // User area 2 1.8V power
      .vssd1(vssd1_core),  // User area 1 digital ground
      .vssd2(vssd2_core),  // User area 2 digital ground	


      // SoC Core Interface
      .porb_h(porb_h),
      .por_l(por_l),
      .rstb_h(rstb_h),
      .clock_core(clock_core),
      .gpio_out_core(gpio_out_core),
      .gpio_in_core(gpio_in_core),
      .gpio_mode0_core(gpio_mode0_core),
      .gpio_mode1_core(gpio_mode1_core),
      .gpio_outenb_core(gpio_outenb_core),
      .gpio_inenb_core(gpio_inenb_core),

      // Flash SPI communication
      .flash_csb_frame(flash_csb_frame),
      .flash_clk_frame(flash_clk_frame),
      .flash_csb_oeb(flash_csb_oeb),
      .flash_clk_oeb(flash_clk_oeb),
      .flash_io0_oeb(flash_io0_oeb),
      .flash_io1_oeb(flash_io1_oeb),
      .flash_io0_ieb(flash_io0_ieb),
      .flash_io1_ieb(flash_io1_ieb),
      .flash_io0_do(flash_io0_do),
      .flash_io1_do(flash_io1_do),
      .flash_io0_di(flash_io0_di),
      .flash_io1_di(flash_io1_di),

      // User project IOs
      .mprj_io_in(mprj_io_in),
      .mprj_io_out(mprj_io_out),
      .mprj_io_oeb(mprj_io_oeb),
      .mprj_io_inp_dis(mprj_io_inp_dis),
      .mprj_io_ib_mode_sel(mprj_io_ib_mode_sel),
      .mprj_io_vtrip_sel(mprj_io_vtrip_sel),
      .mprj_io_slow_sel(mprj_io_slow_sel),
      .mprj_io_holdover(mprj_io_holdover),
      .mprj_io_analog_en(mprj_io_analog_en),
      .mprj_io_analog_sel(mprj_io_analog_sel),
      .mprj_io_analog_pol(mprj_io_analog_pol),
      .mprj_io_dm(mprj_io_dm),

      // Loopbacks to constant value 1 in the 1.8V domain
      .mprj_io_one(mprj_io_one),

      // User project direct access to gpio pad connections for analog
      // (all but the lowest-numbered 7 pads)
      .mprj_analog_io(user_analog_io)
  );

copyright_block copyright_block();
caravel_logo caravel_logo();
caravel_motto caravel_motto();
open_source open_source();
user_id_textblock user_id_textblock();

endmodule
// `default_nettype wire
// SPDX-FileCopyrightText: 2022 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//	http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/*
 * gpio_signal_buffering_alt ---
 *
 * This macro buffers long wires between housekeeping and the GPIO control
 * blocks at the top level of caravan.  The rule of thumb is to limit any
 * single wire length to approximately 1.3mm.  The physical (manhattan)
 * distances and required buffering are as follows:
 *
 * Breakpoints: 1.3, 2.6, 3.9, 5.2, 6.5, 7.8	(mm)
 * # buffers:     1,   2,   3,   4,   5,   6
 *
 * GPIO #    	wire length (mm)	# buffers
 *------------------------------------------------------
 * GPIO 0	0.4			0
 * GPIO 1	0.2			0
 * GPIO 2	0.0			0
 * GPIO 3	0.3			0
 * GPIO 4	0.5			0
 * GPIO 5	0.7			0
 * GPIO 6	1.0			0
 * GPIO 7	1.4			1	
 * GPIO 8	1.6			1
 * GPIO 9	1.8			1
 * GPIO 10	2.1			1
 * GPIO 11	2.3			1
 * GPIO 12	2.5			1
 * GPIO 13	2.7			2	   RHS	
 *-------------------------------------------------------
 * GPIO 25	6.1			4	   LHS
 * GPIO 26	5.9			4
 * GPIO 27	5.7			4
 * GPIO 28	5.5			4
 * GPIO 29	5.3			4
 * GPIO 30	5.1			3
 * GPIO 31	4.8			3
 * GPIO 32	4.2			3
 * GPIO 33	4.0			3
 * GPIO 34	3.8			2
 * GPIO 35	3.5			2
 * GPIO 36	3.3			2
 * GPIO 37	3.4			2
 *------------------------------------------------------
 *	       total number of buffers: 48 (x2 for input and output)
 *
 * OEB lines go to GPIO 0 and 1 (no buffers needed) and GPIO 35-37
 * (2 buffers needed), so OEB lines need 6 additional buffers.
 *
 * The assumption is that all GPIOs on the left-hand side of the chip are
 * routed by taking wires left from the housekeeping across the top of the
 * SoC to the left side, and then up to the destination.  Right-hand side
 * connections go directly up the right side from the housekeeping block.
 *
 * Note that signal names are related to the signal being passed through;
 * "in" and "out" refer to the direction of the signal relative to the
 * housekeeping block in the top level.  For this macro, unbuffered signals
 * "unbuf" are the inputs, and buffered signals "buf" are the outputs.
 */

module gpio_signal_buffering_alt (

    vccd,
    vssd,

    mgmt_io_in_unbuf,
    mgmt_io_out_unbuf,
    mgmt_io_oeb_buf,
    mgmt_io_in_buf,
    mgmt_io_out_buf,
    mgmt_io_oeb_unbuf
);


    input  vccd;
    input  vssd;


    /* NOTE:  To match the indices of the same signals in the
     * top level, add 35 to all OEB lines and add 7 to all in
     * and out lines up to 14, and add 18 to all in and out
     * lines above that.
     */
    input  [19:0] mgmt_io_in_unbuf;
    input  [19:0] mgmt_io_out_unbuf;
    input  [2:0] mgmt_io_oeb_unbuf;
    output [2:0] mgmt_io_oeb_buf;
    output [19:0] mgmt_io_in_buf;
    output [19:0] mgmt_io_out_buf;

    /* Instantiate 48 + 48 + 6 = 101 buffers of size 8 */

    wire [101:0] buf_in;
    wire [101:0] buf_out;

    sky130_fd_sc_hd__buf_8 signal_buffers [101:0] (
        
	    .VPWR(vccd),
	    .VGND(vssd),
	    .VPB(vccd),
	    .VNB(vssd),
	
	.A(buf_in),
	.X(buf_out)
    );

    /* Now chain them all together */

    //----------------------------------------
    // mgmt_io_in, right-hand side
    //----------------------------------------

    assign buf_in[0] = mgmt_io_in_unbuf[0];
    assign mgmt_io_in_buf[0] = buf_out[0];

    assign buf_in[1] = mgmt_io_in_unbuf[1];
    assign mgmt_io_in_buf[1] = buf_out[1];

    assign buf_in[2] = mgmt_io_in_unbuf[2];
    assign mgmt_io_in_buf[2] = buf_out[2];

    assign buf_in[3] = mgmt_io_in_unbuf[3];
    assign mgmt_io_in_buf[3] = buf_out[3];

    assign buf_in[4] = mgmt_io_in_unbuf[4];
    assign mgmt_io_in_buf[4] = buf_out[4];

    assign buf_in[5] = mgmt_io_in_unbuf[5];
    assign mgmt_io_in_buf[5] = buf_out[5];

    assign buf_in[6] = mgmt_io_in_unbuf[6];
    assign buf_in[7] = buf_out[6];
    assign mgmt_io_in_buf[6] = buf_out[7];

    //----------------------------------------
    // mgmt_io_in, left-hand side
    //----------------------------------------

    assign buf_in[8] = mgmt_io_in_unbuf[7];
    assign buf_in[9] = buf_out[8];
    assign buf_in[10] = buf_out[9];
    assign buf_in[11] = buf_out[10];
    assign mgmt_io_in_buf[7] = buf_out[11];

    assign buf_in[12] = mgmt_io_in_unbuf[8];
    assign buf_in[13] = buf_out[12];
    assign buf_in[14] = buf_out[13];
    assign buf_in[15] = buf_out[14];
    assign mgmt_io_in_buf[8] = buf_out[15];

    assign buf_in[16] = mgmt_io_in_unbuf[9];
    assign buf_in[17] = buf_out[16];
    assign buf_in[18] = buf_out[17];
    assign buf_in[19] = buf_out[18];
    assign mgmt_io_in_buf[9] = buf_out[19];

    assign buf_in[20] = mgmt_io_in_unbuf[10];
    assign buf_in[21] = buf_out[20];
    assign buf_in[22] = buf_out[21];
    assign buf_in[23] = buf_out[22];
    assign mgmt_io_in_buf[10] = buf_out[23];

    assign buf_in[24] = mgmt_io_in_unbuf[11];
    assign buf_in[25] = buf_out[24];
    assign buf_in[26] = buf_out[25];
    assign buf_in[27] = buf_out[26];
    assign mgmt_io_in_buf[11] = buf_out[27];

    assign buf_in[28] = mgmt_io_in_unbuf[12];
    assign buf_in[29] = buf_out[28];
    assign buf_in[30] = buf_out[29];
    assign mgmt_io_in_buf[12] = buf_out[30];

    assign buf_in[31] = mgmt_io_in_unbuf[13];
    assign buf_in[32] = buf_out[31];
    assign buf_in[33] = buf_out[32];
    assign mgmt_io_in_buf[13] = buf_out[33];

    assign buf_in[34] = mgmt_io_in_unbuf[14];
    assign buf_in[35] = buf_out[34];
    assign buf_in[36] = buf_out[35];
    assign mgmt_io_in_buf[14] = buf_out[36];

    assign buf_in[37] = mgmt_io_in_unbuf[15];
    assign buf_in[38] = buf_out[37];
    assign buf_in[39] = buf_out[38];
    assign mgmt_io_in_buf[15] = buf_out[39];

    assign buf_in[40] = mgmt_io_in_unbuf[16];
    assign buf_in[41] = buf_out[40];
    assign mgmt_io_in_buf[16] = buf_out[41];

    assign buf_in[42] = mgmt_io_in_unbuf[17];
    assign buf_in[43] = buf_out[42];
    assign mgmt_io_in_buf[17] = buf_out[43];

    assign buf_in[44] = mgmt_io_in_unbuf[18];
    assign buf_in[45] = buf_out[44];
    assign mgmt_io_in_buf[18] = buf_out[45];

    assign buf_in[46] = mgmt_io_in_unbuf[19];
    assign buf_in[47] = buf_out[46];
    assign mgmt_io_in_buf[19] = buf_out[47];

    //----------------------------------------
    // mgmt_io_out, right-hand side
    //----------------------------------------

    assign buf_in[48] = mgmt_io_out_unbuf[0];
    assign mgmt_io_out_buf[0] = buf_out[48];

    assign buf_in[49] = mgmt_io_out_unbuf[1];
    assign mgmt_io_out_buf[1] = buf_out[49];

    assign buf_in[50] = mgmt_io_out_unbuf[2];
    assign mgmt_io_out_buf[2] = buf_out[50];

    assign buf_in[51] = mgmt_io_out_unbuf[3];
    assign mgmt_io_out_buf[3] = buf_out[51];

    assign buf_in[52] = mgmt_io_out_unbuf[4];
    assign mgmt_io_out_buf[4] = buf_out[52];

    assign buf_in[53] = mgmt_io_out_unbuf[5];
    assign mgmt_io_out_buf[5] = buf_out[53];

    assign buf_in[54] = mgmt_io_out_unbuf[6];
    assign buf_in[55] = buf_out[54];
    assign mgmt_io_out_buf[6] = buf_out[55];

    //----------------------------------------
    // mgmt_io_out, left-hand side
    //----------------------------------------

    assign buf_in[56] = mgmt_io_out_unbuf[7];
    assign buf_in[57] = buf_out[56];
    assign buf_in[58] = buf_out[57];
    assign buf_in[59] = buf_out[58];
    assign mgmt_io_out_buf[7] = buf_out[59];

    assign buf_in[60] = mgmt_io_out_unbuf[8];
    assign buf_in[61] = buf_out[60];
    assign buf_in[62] = buf_out[61];
    assign buf_in[63] = buf_out[62];
    assign mgmt_io_out_buf[8] = buf_out[63];

    assign buf_in[64] = mgmt_io_out_unbuf[9];
    assign buf_in[65] = buf_out[64];
    assign buf_in[66] = buf_out[65];
    assign buf_in[67] = buf_out[66];
    assign mgmt_io_out_buf[9] = buf_out[67];

    assign buf_in[68] = mgmt_io_out_unbuf[10];
    assign buf_in[69] = buf_out[68];
    assign buf_in[70] = buf_out[69];
    assign buf_in[71] = buf_out[70];
    assign mgmt_io_out_buf[10] = buf_out[71];

    assign buf_in[72] = mgmt_io_out_unbuf[11];
    assign buf_in[73] = buf_out[72];
    assign buf_in[74] = buf_out[73];
    assign buf_in[75] = buf_out[74];
    assign mgmt_io_out_buf[11] = buf_out[75];

    assign buf_in[76] = mgmt_io_out_unbuf[12];
    assign buf_in[77] = buf_out[76];
    assign buf_in[78] = buf_out[77];
    assign mgmt_io_out_buf[12] = buf_out[78];

    assign buf_in[79] = mgmt_io_out_unbuf[13];
    assign buf_in[80] = buf_out[79];
    assign buf_in[81] = buf_out[80];
    assign mgmt_io_out_buf[13] = buf_out[81];

    assign buf_in[82] = mgmt_io_out_unbuf[14];
    assign buf_in[83] = buf_out[82];
    assign buf_in[84] = buf_out[83];
    assign mgmt_io_out_buf[14] = buf_out[84];

    assign buf_in[85] = mgmt_io_out_unbuf[15];
    assign buf_in[86] = buf_out[85];
    assign buf_in[87] = buf_out[86];
    assign mgmt_io_out_buf[15] = buf_out[87];

    assign buf_in[88] = mgmt_io_out_unbuf[16];
    assign buf_in[89] = buf_out[88];
    assign mgmt_io_out_buf[16] = buf_out[89];

    assign buf_in[90] = mgmt_io_out_unbuf[17];
    assign buf_in[91] = buf_out[90];
    assign mgmt_io_out_buf[17] = buf_out[91];

    assign buf_in[92] = mgmt_io_out_unbuf[18];
    assign buf_in[93] = buf_out[92];
    assign mgmt_io_out_buf[18] = buf_out[93];

    assign buf_in[94] = mgmt_io_out_unbuf[19];
    assign buf_in[95] = buf_out[94];
    assign mgmt_io_out_buf[19] = buf_out[95];

    //----------------------------------------
    // mgmt_io_oeb, left-hand side (only)
    //----------------------------------------

    assign buf_in[96] = mgmt_io_oeb_unbuf[0];
    assign buf_in[97] = buf_out[96];
    assign mgmt_io_oeb_buf[0] = buf_out[97];

    assign buf_in[98] = mgmt_io_oeb_unbuf[1];
    assign buf_in[99] = buf_out[98];
    assign mgmt_io_oeb_buf[1] = buf_out[99];

    assign buf_in[100] = mgmt_io_oeb_unbuf[2];
    assign buf_in[101] = buf_out[100];
    assign mgmt_io_oeb_buf[2] = buf_out[101];

    sky130_ef_sc_hd__decap_12 sigbuf_decaps [59:0] (
    
        .VPWR(vccd),
        .VGND(vssd),
        .VPB(vccd),
        .VNB(vssd)
    
    );

endmodule
// `default_nettype none
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0
/*--------------------------------------------------------------*/
/* caravan, a project harness for the Google/SkyWater sky130	*/
/* fabrication process and open source PDK.  caravan is an 	*/
/* alternative architecture to caravel that has simple straight	*/
/* through connections replacing the GPIO pads on the top side	*/
/* of the padframe.  A total of 11 pads are converted from GPIO	*/
/* to analog, leaving 27 GPIO.					*/
/*                                                          	*/
/* Copyright 2021 efabless, Inc.                            	*/
/* Written by Tim Edwards, December 2019                    	*/
/* and Mohamed Shalan, August 2020			    	*/
/* This file is open source hardware released under the     	*/
/* Apache 2.0 license.  See file LICENSE.                   	*/
/*                                                          	*/
/*--------------------------------------------------------------*/

/*--------------------------------------------------------------*/
/* Derived types for the array bounds on the two digital and	*/
/* two analog pad arrays.  As defined above, the sections have	*/
/* the number of pads as follows:				*/
/*								*/
/*	DIG2 : 13 GPIO pads					*/
/*	ANA2 : 6  analog pads					*/
/*	ANA1 : 5  analog pads					*/
/*	DIG1 : 14 GPIO pads					*/
/*								*/
/* This makes a total of 38 pads = `MPRJ_IO_PADS		*/
/* The pads are still designated as mprj_io[37:0] around the	*/
/* padframe.  The SoC core remains the same, so the programming	*/
/* of the digital signals remains the same, but the values for	*/
/* GPIO 14-24 (indexed from 0) are not used.			*/
/*--------------------------------------------------------------*/












/*--------------------------------------------------------------*/
/*--------------------------------------------------------------*/

module caravan (
    
        inout vddio,	// Common 3.3V padframe/ESD power
        inout vddio_2,	// Common 3.3V padframe/ESD power
        inout vssio,	// Common padframe/ESD ground
        inout vssio_2,	// Common padframe/ESD ground
        inout vdda,		// Management 3.3V power
        inout vssa,		// Common analog ground
        inout vccd,		// Management/Common 1.8V power
        inout vssd,		// Common digital ground
        inout vdda1,	// User area 1 3.3V power
        inout vdda1_2,	// User area 1 3.3V power
        inout vdda2,	// User area 2 3.3V power
        inout vssa1,	// User area 1 analog ground
        inout vssa1_2,	// User area 1 analog ground
        inout vssa2,	// User area 2 analog ground
        inout vccd1,	// User area 1 1.8V power
        inout vccd2,	// User area 2 1.8V power
        inout vssd1,	// User area 1 digital ground
        inout vssd2,	// User area 2 digital ground
    

    inout gpio,			// Used for external LDO control
    inout [(19 + 19)-1:0] mprj_io,
    input clock,	    	// CMOS core clock input, not a crystal
    input resetb,

    // Note that only two pins are available on the flash so dual and
    // quad flash modes are not available.

    output flash_csb,
    output flash_clk,
    output flash_io0,
    output flash_io1
);

    //------------------------------------------------------------
    // This value is uniquely defined for each user project.
    //------------------------------------------------------------
    parameter USER_PROJECT_ID = 32'h00000000;

    /*
     *---------------------------------------------------------------------
     * These pins are overlaid on mprj_io space.  They have the function
     * below when the management processor is in reset, or in the default
     * configuration.  They are assigned to uses in the user space by the
     * configuration program running off of the SPI flash.  Note that even
     * when the user has taken control of these pins, they can be restored
     * to the original use by setting the resetb pin low.  The SPI pins and
     * UART pins can be connected directly to an FTDI chip as long as the
     * FTDI chip sets these lines to high impedence (input function) at
     * all times except when holding the chip in reset.
     *
     * JTAG      = mprj_io[0]		(inout)
     * SDO 	 = mprj_io[1]		(output)
     * SDI 	 = mprj_io[2]		(input)
     * CSB 	 = mprj_io[3]		(input)
     * SCK	 = mprj_io[4]		(input)
     * ser_rx    = mprj_io[5]		(input)
     * ser_tx    = mprj_io[6]		(output)
     * irq 	 = mprj_io[7]		(input)
     *
     * spi_sck    = mprj_io[32]         (output)
     * spi_csb    = mprj_io[33]         (output)
     * spi_sdi    = mprj_io[34]         (input)
     * spi_sdo    = mprj_io[35]         (output)
     * flash_io2  = mprj_io[36]         (inout)
     * flash_io3  = mprj_io[37]         (inout)
     *
     * These pins are reserved for any project that wants to incorporate
     * its own processor and flash controller.  While a user project can
     * technically use any available I/O pins for the purpose, these
     * four pins connect to a pass-through mode from the SPI slave (pins
     * 1-4 above) so that any SPI flash connected to these specific pins
     * can be accessed through the SPI slave even when the processor is in
     * reset.
     *
     * user_flash_csb = mprj_io[8]
     * user_flash_sck = mprj_io[9]
     * user_flash_io0 = mprj_io[10]
     * user_flash_io1 = mprj_io[11]
     *
     *---------------------------------------------------------------------
     */

    // One-bit GPIO dedicated to management SoC (outside of user control)
    wire gpio_out_core;
    wire gpio_in_core;
    wire gpio_mode0_core;
    wire gpio_mode1_core;
    wire gpio_outenb_core;
    wire gpio_inenb_core;

    // 27 GPIO pads with full controls
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_inp_dis;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_oeb;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_ib_mode_sel;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_vtrip_sel;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_slow_sel;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_holdover;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_analog_en;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_analog_sel;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_analog_pol;
    wire [((19 + 19)-(5 + 6))*3-1:0] mprj_io_dm;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_in;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_in_3v3;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_out;
    wire [(19 + 19)-(5 + 6)-1:0] mprj_io_one;
    wire [7:0] mprj_io_zero;

    // User Project Control (user-facing)
    // 27 GPIO bidirectional with in/out/oeb and a 3.3V copy of the input
    wire [(19 + 19)-(5 + 6)-1:0] user_io_oeb;
    wire [(19 + 19)-(5 + 6)-1:0] user_io_in;
    wire [(19 + 19)-(5 + 6)-1:0] user_io_out;
    wire [(19 + 19)-(5 + 6)-1:0] user_io_in_3v3;

    // 18 direct connections to GPIO for low-frequency, low-voltage analog
    wire [(19 + 19)-(5 + 6)-10:0] user_gpio_analog;
    wire [(19 + 19)-(5 + 6)-10:0] user_gpio_noesd;

    // 3 power supply ESD clamps for user applications
    wire [2:0] user_clamp_high;
    wire [2:0] user_clamp_low;

    // 11 core connections to the analog pads
    wire [(5 + 6)-1:0] user_analog;

    /* Padframe control signals */
    wire [19-5-1:0] gpio_serial_link_1;
    wire [19-6-1:0] gpio_serial_link_2;
    wire mprj_io_loader_resetn;
    wire mprj_io_loader_clock;
    wire mprj_io_loader_strobe;
    wire mprj_io_loader_data_1;		/* user1 side serial loader */
    wire mprj_io_loader_data_2;		/* user2 side serial loader */

    // User Project Control management I/O
    // There are two types of GPIO connections:
    // (1) Full Bidirectional: Management connects to in, out, and oeb
    //     Uses:  JTAG and SDO
    // (2) Selectable bidirectional:  Management connects to in and out,
    //	   which are tied together.  oeb is grounded (oeb from the
    //	   configuration is used)

    // SDI 	 = mprj_io[2]		(input)
    // CSB 	 = mprj_io[3]		(input)
    // SCK	 = mprj_io[4]		(input)
    // ser_rx    = mprj_io[5]		(input)
    // ser_tx    = mprj_io[6]		(output)
    // irq 	 = mprj_io[7]		(input)

    wire [(19 + 19)-1:0] mgmt_io_in;	/* two- and three-pin data in */
    wire [(19 + 19)-1:0] mgmt_io_out;	/* two- and three-pin data out */
    wire [(19 + 19)-1:0] mgmt_io_oeb;	/* output enable, used only by	*/
						/* three-pin interfaces		*/
    wire [(2 + 2)-1:0] pwr_ctrl_nc;	/* no-connects */

    /* Buffers are placed between housekeeping and gpio_control_block		*/
    /* instances to mitigate timing issues on very long (> 1.5mm) wires.	*/
    wire [(19 + 19)-1:0] mgmt_io_in_hk;	/* mgmt_io_in at housekeeping	*/
    wire [(19 + 19)-1:0] mgmt_io_out_hk;	/* mgmt_io_out at housekeeping	*/
    wire [(19 + 19)-1:0] mgmt_io_oeb_hk;	/* mgmt_io_oeb at housekeeping	*/

    wire clock_core;

    // Power-on-reset signal.  The reset pad generates the sense-inverted
    // reset at 3.3V.  The 1.8V signal and the inverted 1.8V signal are
    // derived.

    wire porb_h;
    wire porb_l;
    wire por_l;

    wire rstb_h;
    wire rstb_l;

    // Flash SPI communication (managment SoC to housekeeping)
    wire flash_clk_core,     flash_csb_core;
    wire flash_clk_oeb_core, flash_csb_oeb_core;
    wire flash_io0_oeb_core, flash_io1_oeb_core;
    wire flash_io2_oeb_core, flash_io3_oeb_core;
    wire flash_io0_ieb_core, flash_io1_ieb_core;
    wire flash_io2_ieb_core, flash_io3_ieb_core;
    wire flash_io0_do_core,  flash_io1_do_core;
    wire flash_io2_do_core,  flash_io3_do_core;
    wire flash_io0_di_core,  flash_io1_di_core;
    wire flash_io2_di_core,  flash_io3_di_core;

    // Flash SPI communication
    wire flash_clk_frame;
    wire flash_csb_frame;
    wire flash_clk_oeb, flash_csb_oeb;
    wire flash_io0_oeb, flash_io1_oeb;
    wire flash_io0_ieb, flash_io1_ieb;
    wire flash_io0_do,  flash_io1_do;
    wire flash_io0_di,  flash_io1_di;

	// Flash buffered signals
    wire flash_clk_frame_buf;
    wire flash_csb_frame_buf;
    wire flash_io0_oeb_buf, flash_io1_oeb_buf;
    wire flash_io0_ieb_buf, flash_io1_ieb_buf;
    wire flash_io0_do_buf,  flash_io1_do_buf;
    wire flash_io0_di_buf,  flash_io1_di_buf;

	// Clock and reset buffered signals
	wire caravel_clk_buf;
	wire caravel_rstn_buf;
	wire clock_core_buf;

	// SoC pass through buffered signals
	wire mprj_io_loader_clock_buf;
	wire mprj_io_loader_strobe_buf;
	wire mprj_io_loader_resetn_buf;
	wire mprj_io_loader_data_2_buf;
	wire rstb_l_buf;
	wire por_l_buf;
	wire porb_h_buf;

    // SoC core
    wire caravel_clk;
    wire caravel_clk2;
    wire caravel_rstn;
	
	// top-level buffers
	buff_flash_clkrst flash_clkrst_buffers (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	
	.in_n({
		caravel_clk,
		caravel_rstn,
		flash_clk_frame, 
		flash_csb_frame, 
		flash_clk_oeb, 
		flash_csb_oeb, 
		flash_io0_oeb, 
		flash_io1_oeb,
		flash_io0_ieb, 
		flash_io1_ieb,
		flash_io0_do,  
		flash_io1_do }), 
	.in_s({
		clock_core,
		flash_io1_di, 
		flash_io0_di }),
	.out_s({ 
		caravel_clk_buf,
		caravel_rstn_buf,
		flash_clk_frame_buf, 
		flash_csb_frame_buf, 
		flash_clk_oeb_buf, 
		flash_csb_oeb_buf, 
		flash_io0_oeb_buf, 
		flash_io1_oeb_buf,
		flash_io0_ieb_buf, 
		flash_io1_ieb_buf,
		flash_io0_do_buf,  
		flash_io1_do_buf }), 
	.out_n({
		clock_core_buf,
		flash_io1_di_buf, 
		flash_io0_di_buf })
	);







    assign mgmt_io_in_hk[6:0] = mgmt_io_in[6:0];
    assign mgmt_io_out[6:0] = mgmt_io_out_hk[6:0];
    assign mgmt_io_oeb[34:0] = mgmt_io_oeb_hk[34:0];

    /* The following are tied to ground through the zero value	*/
    /* outputs of the closest GPIO control blocks.  Tie two 	*/
    /* inputs to one zero value output so that the wires from	*/
    /* the GPIOs to housekeeping don't get too long.		*/
    assign mgmt_io_in_hk[24:14] = {mprj_io_zero[5],
		mprj_io_zero[4], mprj_io_zero[4],
		mprj_io_zero[3], mprj_io_zero[3],
		mprj_io_zero[2], mprj_io_zero[2],
		mprj_io_zero[1], mprj_io_zero[1],
		mprj_io_zero[0], mprj_io_zero[0]};

    /* The following are no-connects in caravan (no associated GPIO) */
    assign mgmt_io_out[24:14] = mgmt_io_out_hk[24:14];

    gpio_signal_buffering_alt sigbuf (
	
	    .vccd(vccd_core),
	    .vssd(vssd_core),
	
	.mgmt_io_in_unbuf({mgmt_io_in[37:25],mgmt_io_in[13:7]}),
	.mgmt_io_out_unbuf({mgmt_io_out_hk[37:25],mgmt_io_out_hk[13:7]}),
	.mgmt_io_oeb_unbuf(mgmt_io_oeb_hk[37:35]),
	.mgmt_io_in_buf({mgmt_io_in_hk[37:25],mgmt_io_in_hk[13:7]}),
	.mgmt_io_out_buf({mgmt_io_out[37:25],mgmt_io_out[13:7]}),
	.mgmt_io_oeb_buf(mgmt_io_oeb[37:35])
    );


    chip_io_alt #(
	.ANALOG_PADS_1(5),
	.ANALOG_PADS_2(6)
    ) padframe (
	
		// Package Pins
		.vddio_pad	(vddio),		// Common padframe/ESD supply
		.vddio_pad2	(vddio_2),
		.vssio_pad	(vssio),		// Common padframe/ESD ground
		.vssio_pad2	(vssio_2),
		.vccd_pad	(vccd),			// Common 1.8V supply
		.vssd_pad	(vssd),			// Common digital ground
		.vdda_pad	(vdda),			// Management analog 3.3V supply
		.vssa_pad	(vssa),			// Management analog ground
		.vdda1_pad	(vdda1),		// User area 1 3.3V supply
		.vdda1_pad2	(vdda1_2),		
		.vdda2_pad	(vdda2),		// User area 2 3.3V supply
		.vssa1_pad	(vssa1),		// User area 1 analog ground
		.vssa1_pad2	(vssa1_2),
		.vssa2_pad	(vssa2),		// User area 2 analog ground
		.vccd1_pad	(vccd1),		// User area 1 1.8V supply
		.vccd2_pad	(vccd2),		// User area 2 1.8V supply
		.vssd1_pad	(vssd1),		// User area 1 digital ground
		.vssd2_pad	(vssd2),		// User area 2 digital ground
        .vddio	(vddio_core),
        .vssio	(vssio_core),
        .vdda	(vdda_core),
        .vssa	(vssa_core),
        .vccd	(vccd_core),
        .vssd	(vssd_core),
        .vdda1	(vdda1_core),
        .vdda2	(vdda2_core),
        .vssa1	(vssa1_core),
        .vssa2	(vssa2_core),
        .vccd1	(vccd1_core),
        .vccd2	(vccd2_core),
        .vssd1	(vssd1_core),
        .vssd2	(vssd2_core),
	
	
	// Core Side Pins
	.gpio(gpio),
	.mprj_io(mprj_io),
	.clock(clock),
	.resetb(resetb),
	.flash_csb(flash_csb),
	.flash_clk(flash_clk),
	.flash_io0(flash_io0),
	.flash_io1(flash_io1),
	// SoC Core Interface
	.porb_h(porb_h),
	.por(por_l_buf),
	.resetb_core_h(rstb_h),
	.clock_core(clock_core),
	.gpio_out_core(gpio_out_core),
	.gpio_in_core(gpio_in_core),
	.gpio_mode0_core(gpio_mode0_core),
	.gpio_mode1_core(gpio_mode1_core),
	.gpio_outenb_core(gpio_outenb_core),
	.gpio_inenb_core(gpio_inenb_core),
	.flash_csb_core(flash_csb_frame_buf),
	.flash_clk_core(flash_clk_frame_buf),
	.flash_csb_oeb_core(flash_csb_oeb_buf),
	.flash_clk_oeb_core(flash_clk_oeb_buf),
	.flash_io0_oeb_core(flash_io0_oeb_buf),
	.flash_io1_oeb_core(flash_io1_oeb_buf),
	.flash_io0_ieb_core(flash_io0_ieb_buf),
	.flash_io1_ieb_core(flash_io1_ieb_buf),
	.flash_io0_do_core(flash_io0_do_buf),
	.flash_io1_do_core(flash_io1_do_buf),
	.flash_io0_di_core(flash_io0_di),
	.flash_io1_di_core(flash_io1_di),
	.mprj_io_one(mprj_io_one),
	.mprj_io_in(mprj_io_in),
	.mprj_io_in_3v3(mprj_io_in_3v3),
	.mprj_io_out(mprj_io_out),
	.mprj_io_oeb(mprj_io_oeb),
	.mprj_io_inp_dis(mprj_io_inp_dis),
	.mprj_io_ib_mode_sel(mprj_io_ib_mode_sel),
	.mprj_io_vtrip_sel(mprj_io_vtrip_sel),
	.mprj_io_slow_sel(mprj_io_slow_sel),
	.mprj_io_holdover(mprj_io_holdover),
	.mprj_io_analog_en(mprj_io_analog_en),
	.mprj_io_analog_sel(mprj_io_analog_sel),
	.mprj_io_analog_pol(mprj_io_analog_pol),
	.mprj_io_dm(mprj_io_dm),
	.mprj_gpio_analog(user_gpio_analog),
	.mprj_gpio_noesd(user_gpio_noesd),
	.mprj_analog(user_analog),
	.mprj_clamp_high(user_clamp_high),
	.mprj_clamp_low(user_clamp_low)
    );



    wire [7:0] spi_ro_config_core;

    // LA signals
    wire [127:0] la_data_in_user;  // From CPU to MPRJ
    wire [127:0] la_data_in_mprj;  // From MPRJ to CPU
    wire [127:0] la_data_out_mprj; // From CPU to MPRJ
    wire [127:0] la_data_out_user; // From MPRJ to CPU
    wire [127:0] la_oenb_user;     // From CPU to MPRJ
    wire [127:0] la_oenb_mprj;	   // From CPU to MPRJ
    wire [127:0] la_iena_mprj;     // From CPU only

    wire [2:0]   user_irq;	   // From MPRJ to CPU
    wire [2:0]   user_irq_core;
    wire [2:0]   user_irq_ena;
    wire [2:0]	 irq_spi;	   // From SPI and external pins

    // Exported Wishbone Bus (processor facing)
    wire mprj_iena_wb;
    wire mprj_cyc_o_core;
    wire mprj_stb_o_core;
    wire mprj_we_o_core;
    wire [3:0] mprj_sel_o_core;
    wire [31:0] mprj_adr_o_core;
    wire [31:0] mprj_dat_o_core;
    wire 	mprj_ack_i_core;
    wire [31:0] mprj_dat_i_core;

    wire [31:0] hk_dat_i;
    wire hk_ack_i;
    wire hk_stb_o;
    wire hk_cyc_o;

    // Exported Wishbone Bus (user area facing)
    wire 	mprj_cyc_o_user;
    wire 	mprj_stb_o_user;
    wire 	mprj_we_o_user;
    wire [3:0]  mprj_sel_o_user;
    wire [31:0] mprj_adr_o_user;
    wire [31:0] mprj_dat_o_user;
    wire [31:0]	mprj_dat_i_user;
    wire 	mprj_ack_i_user;

    // Mask revision
    wire [31:0] mask_rev;

    wire 	mprj_clock;
    wire 	mprj_clock2;
    wire 	mprj_reset;

    // Power monitoring
    wire	mprj_vcc_pwrgood;
    wire	mprj2_vcc_pwrgood;
    wire	mprj_vdd_pwrgood;
    wire	mprj2_vdd_pwrgood;









    // Management processor (wrapper).  Any management core
    // implementation must match this pinout.

    // Pass thru clock and reset
    wire 	clk_passthru;
    wire 	resetn_passthru;

    // NC passthru signal porb_h
    wire porb_h_out_nc;

    mgmt_core_wrapper soc (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	

	// SoC pass through buffered signals
	.serial_clock_in(mprj_io_loader_clock),
	.serial_clock_out(mprj_io_loader_clock_buf),
	.serial_load_in(mprj_io_loader_strobe),
	.serial_load_out(mprj_io_loader_strobe_buf),
	.serial_resetn_in(mprj_io_loader_resetn),
	.serial_resetn_out(mprj_io_loader_resetn_buf),
	.serial_data_2_in(mprj_io_loader_data_2),
	.serial_data_2_out(mprj_io_loader_data_2_buf),
	.rstb_l_in(rstb_l),
	.rstb_l_out(rstb_l_buf),
	.porb_h_in(por_l),		// NOTE: purposefully tied off to por_l_in
	.porb_h_out(porb_h_out_nc),
	.por_l_in(por_l),
	.por_l_out(por_l_buf),

	// Clock and reset
	.core_clk(caravel_clk_buf),
	.core_rstn(caravel_rstn_buf),

    // Pass thru Clock and reset
	.clk_in(caravel_clk_buf),
	.resetn_in(caravel_rstn_buf),
	.clk_out(clk_passthru),
	.resetn_out(resetn_passthru),

	// GPIO (1 pin)
	.gpio_out_pad(gpio_out_core),
	.gpio_in_pad(gpio_in_core),
	.gpio_mode0_pad(gpio_mode0_core),
	.gpio_mode1_pad(gpio_mode1_core),
	.gpio_outenb_pad(gpio_outenb_core),
	.gpio_inenb_pad(gpio_inenb_core),

	// Primary SPI flash controller
	.flash_csb(flash_csb_core),
	.flash_clk(flash_clk_core),
	.flash_io0_oeb(flash_io0_oeb_core),
	.flash_io0_di(flash_io0_di_core),
	.flash_io0_do(flash_io0_do_core),
	.flash_io1_oeb(flash_io1_oeb_core),
	.flash_io1_di(flash_io1_di_core),
	.flash_io1_do(flash_io1_do_core),
	.flash_io2_oeb(flash_io2_oeb_core),
	.flash_io2_di(flash_io2_di_core),
	.flash_io2_do(flash_io2_do_core),
	.flash_io3_oeb(flash_io3_oeb_core),
	.flash_io3_di(flash_io3_di_core),
	.flash_io3_do(flash_io3_do_core),

	// Exported Wishbone Bus
	.mprj_wb_iena(mprj_iena_wb),
	.mprj_cyc_o(mprj_cyc_o_core),
	.mprj_stb_o(mprj_stb_o_core),
	.mprj_we_o(mprj_we_o_core),
	.mprj_sel_o(mprj_sel_o_core),
	.mprj_adr_o(mprj_adr_o_core),
	.mprj_dat_o(mprj_dat_o_core),
	.mprj_ack_i(mprj_ack_i_core),
	.mprj_dat_i(mprj_dat_i_core),

	.hk_stb_o(hk_stb_o),
	.hk_cyc_o(hk_cyc_o),
	.hk_dat_i(hk_dat_i),
	.hk_ack_i(hk_ack_i),

	// IRQ
	.irq({irq_spi, user_irq}),
	.user_irq_ena(user_irq_ena),

	// Module status (these may or may not be implemented)
	.qspi_enabled(qspi_enabled),
	.uart_enabled(uart_enabled),
	.spi_enabled(spi_enabled),
	.debug_mode(debug_mode),

	// Module I/O (these may or may not be implemented)
	// UART
	.ser_tx(ser_tx),
	.ser_rx(ser_rx),
	// SPI master
	.spi_sdi(spi_sdi),
	.spi_csb(spi_csb),
	.spi_sck(spi_sck),
	.spi_sdo(spi_sdo),
	.spi_sdoenb(spi_sdoenb),
	// Debug
	.debug_in(debug_in),
	.debug_out(debug_out),
	.debug_oeb(debug_oeb),
	// Logic analyzer
	.la_input(la_data_in_mprj),
	.la_output(la_data_out_mprj),
	.la_oenb(la_oenb_mprj),
	.la_iena(la_iena_mprj),









	// Trap status
	.trap(trap)
    );

    /* Clock and reset to user space are passed through a tristate	*/
    /* buffer like the above, but since they are intended to be		*/
    /* always active, connect the enable to the logic-1 output from	*/
    /* the vccd1 domain.						*/

    mgmt_protect mgmt_buffers (
	
	    .vccd(vccd_core),
	    .vssd(vssd_core),
	    .vccd1(vccd1_core),
	    .vssd1(vssd1_core),
	    .vccd2(vccd2_core),
	    .vssd2(vssd2_core),
	    .vdda1(vdda1_core),
	    .vssa1(vssa1_core),
	    .vdda2(vdda2_core),
	    .vssa2(vssa2_core),
	
	.caravel_clk(clk_passthru),
	.caravel_clk2(caravel_clk2),
	.caravel_rstn(resetn_passthru),
	.mprj_iena_wb(mprj_iena_wb),
	.mprj_cyc_o_core(mprj_cyc_o_core),
	.mprj_stb_o_core(mprj_stb_o_core),
	.mprj_we_o_core(mprj_we_o_core),
	.mprj_sel_o_core(mprj_sel_o_core),
	.mprj_adr_o_core(mprj_adr_o_core),
	.mprj_dat_o_core(mprj_dat_o_core),
	.mprj_ack_i_core(mprj_ack_i_core),
	.mprj_dat_i_core(mprj_dat_i_core),
	.user_irq_core(user_irq_core),
	.user_irq_ena(user_irq_ena),
	.la_data_out_core(la_data_out_user),
	.la_data_out_mprj(la_data_out_mprj),
	.la_data_in_core(la_data_in_user),
	.la_data_in_mprj(la_data_in_mprj),
	.la_oenb_mprj(la_oenb_mprj),
	.la_oenb_core(la_oenb_user),
	.la_iena_mprj(la_iena_mprj),

	.user_clock(mprj_clock),
	.user_clock2(mprj_clock2),
	.user_reset(mprj_reset),
	.mprj_cyc_o_user(mprj_cyc_o_user),
	.mprj_stb_o_user(mprj_stb_o_user),
	.mprj_we_o_user(mprj_we_o_user),
	.mprj_sel_o_user(mprj_sel_o_user),
	.mprj_adr_o_user(mprj_adr_o_user),
	.mprj_dat_o_user(mprj_dat_o_user),
	.mprj_dat_i_user(mprj_dat_i_user),
	.mprj_ack_i_user(mprj_ack_i_user),
	.user_irq(user_irq),
	.user1_vcc_powergood(mprj_vcc_pwrgood),
	.user2_vcc_powergood(mprj2_vcc_pwrgood),
	.user1_vdd_powergood(mprj_vdd_pwrgood),
	.user2_vdd_powergood(mprj2_vdd_pwrgood)
    );


    /*--------------------------------------------------*/
    /* Wrapper module around the user project 		*/
    /*--------------------------------------------------*/

    assign user_io_in_3v3 = mprj_io_in_3v3;
	
    user_analog_project_wrapper mprj ( 
	
	     .vdda1(vdda1_core),	// User area 1 3.3V power
	     .vdda2(vdda2_core),	// User area 2 3.3V power
	     .vssa1(vssa1_core),	// User area 1 analog ground
	     .vssa2(vssa2_core),	// User area 2 analog ground
	     .vccd1(vccd1_core),	// User area 1 1.8V power
	     .vccd2(vccd2_core),	// User area 2 1.8V power
	     .vssd1(vssd1_core),	// User area 1 digital ground
	     .vssd2(vssd2_core),	// User area 2 digital ground
	

    	.wb_clk_i(mprj_clock),
    	.wb_rst_i(mprj_reset),

	// MGMT SoC Wishbone Slave
	.wbs_cyc_i(mprj_cyc_o_user),
	.wbs_stb_i(mprj_stb_o_user),
	.wbs_we_i(mprj_we_o_user),
	.wbs_sel_i(mprj_sel_o_user),
	.wbs_adr_i(mprj_adr_o_user),
	.wbs_dat_i(mprj_dat_o_user),
	.wbs_ack_o(mprj_ack_i_user),
	.wbs_dat_o(mprj_dat_i_user),

	// GPIO pad 3-pin interface (plus analog)
	.io_in (user_io_in),
	.io_in_3v3 (user_io_in_3v3),
    	.io_out(user_io_out),
    	.io_oeb(user_io_oeb),
    
        .io_analog(user_analog),
        .io_clamp_high(user_clamp_high),
        .io_clamp_low(user_clamp_low),
    
	.gpio_analog(user_gpio_analog),
	.gpio_noesd(user_gpio_noesd),

	// Logic Analyzer
	.la_data_in(la_data_in_user),
	.la_data_out(la_data_out_user),
	.la_oenb(la_oenb_user),

	// User-accessible power supply clamps

	// Independent clock
	.user_clock2(mprj_clock2),

	// IRQ
	.user_irq(user_irq_core)
    );

    /*--------------------------------------*/
    /* End user project instantiation	*/
    /*--------------------------------------*/

    wire [19-5-1:0] gpio_serial_link_1_shifted;
    wire [19-6-1:0] gpio_serial_link_2_shifted;

    assign gpio_serial_link_1_shifted = {gpio_serial_link_1[19
					-5-2:0],
					 mprj_io_loader_data_1};
    // Note that serial_link_2 is backwards compared to serial_link_1, so it
    // shifts in the other direction.
    assign gpio_serial_link_2_shifted = {mprj_io_loader_data_2_buf,
					 gpio_serial_link_2[19
					-6-1:1]};

    // Propagating clock and reset to mitigate timing and fanout issues
    wire [19-1:0] gpio_clock_1;
    wire [19-1:0] gpio_clock_2;
    wire [19-1:0] gpio_resetn_1;
    wire [19-1:0] gpio_resetn_2;
    wire [19-1:0] gpio_load_1;
    wire [19-1:0] gpio_load_2;
    wire [19-6:0] gpio_clock_1_shifted;
    wire [19-7:0] gpio_clock_2_shifted;
    wire [19-6:0] gpio_resetn_1_shifted;
    wire [19-7:0] gpio_resetn_2_shifted;
    wire [19-6:0] gpio_load_1_shifted;
    wire [19-7:0] gpio_load_2_shifted;

    assign gpio_clock_1_shifted = {gpio_clock_1[19-5-2:0],
				mprj_io_loader_clock};
    assign gpio_clock_2_shifted = {mprj_io_loader_clock_buf,
				gpio_clock_2[19-6-1:1]};
    assign gpio_resetn_1_shifted = {gpio_resetn_1[19-5-2:0],
				mprj_io_loader_resetn};
    assign gpio_resetn_2_shifted = {mprj_io_loader_resetn_buf,
				gpio_resetn_2[19-6-1:1]};
    assign gpio_load_1_shifted = {gpio_load_1[19-5-2:0],
				mprj_io_loader_strobe};
    assign gpio_load_2_shifted = {mprj_io_loader_strobe_buf,
				gpio_load_2[19-6-1:1]};

    wire [2:0] spi_pll_sel;
    wire [2:0] spi_pll90_sel;
    wire [4:0] spi_pll_div;
    wire [25:0] spi_pll_trim;

    // Clocking control

    caravel_clocking clock_ctrl (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	
	.ext_clk_sel(ext_clk_sel),
	.ext_clk(clock_core_buf),
	.pll_clk(pll_clk),
	.pll_clk90(pll_clk90),
	.resetb(rstb_l_buf),
	.sel(spi_pll_sel),
	.sel2(spi_pll90_sel),
	.ext_reset(ext_reset),  // From housekeeping SPI
	.core_clk(caravel_clk),
	.user_clk(caravel_clk2),
	.resetb_sync(caravel_rstn)
    );

    // DCO/Digital Locked Loop

    digital_pll pll (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	
	.resetb(rstb_l_buf),
	.enable(spi_pll_ena),
	.osc(clock_core_buf),
	.clockp({pll_clk, pll_clk90}),
	.div(spi_pll_div),
	.dco(spi_pll_dco_ena),
	.ext_trim(spi_pll_trim)
    );

    // Housekeeping interface

    housekeeping housekeeping (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	

	.wb_clk_i(caravel_clk),
	.wb_rstn_i(caravel_rstn),

	.wb_adr_i(mprj_adr_o_core),
	.wb_dat_i(mprj_dat_o_core),
	.wb_sel_i(mprj_sel_o_core),
	.wb_we_i(mprj_we_o_core),
	.wb_cyc_i(hk_cyc_o),
	.wb_stb_i(hk_stb_o),
	.wb_ack_o(hk_ack_i),
	.wb_dat_o(hk_dat_i),

	.porb(porb_l),

	.pll_ena(spi_pll_ena),
	.pll_dco_ena(spi_pll_dco_ena),
	.pll_div(spi_pll_div),
	.pll_sel(spi_pll_sel),
	.pll90_sel(spi_pll90_sel),
	.pll_trim(spi_pll_trim),
	.pll_bypass(ext_clk_sel),

	.qspi_enabled(qspi_enabled),
	.uart_enabled(uart_enabled),
	.spi_enabled(spi_enabled),
	.debug_mode(debug_mode),

	.ser_tx(ser_tx),
	.ser_rx(ser_rx),

	.spi_sdi(spi_sdi),
	.spi_csb(spi_csb),
	.spi_sck(spi_sck),
	.spi_sdo(spi_sdo),
	.spi_sdoenb(spi_sdoenb),

	.debug_in(debug_in),
	.debug_out(debug_out),
	.debug_oeb(debug_oeb),

	.irq(irq_spi),
	.reset(ext_reset),

	.serial_clock(mprj_io_loader_clock),
	.serial_load(mprj_io_loader_strobe),
	.serial_resetn(mprj_io_loader_resetn),
	.serial_data_1(mprj_io_loader_data_1),
	.serial_data_2(mprj_io_loader_data_2),

	.mgmt_gpio_in(mgmt_io_in_hk),
	.mgmt_gpio_out(mgmt_io_out_hk),
	.mgmt_gpio_oeb(mgmt_io_oeb_hk),

	.pwr_ctrl_out(pwr_ctrl_nc),        /* Not used in this version */

	.trap(trap),

	.user_clock(caravel_clk2),

	.mask_rev_in(mask_rev),

	.spimemio_flash_csb(flash_csb_core),
	.spimemio_flash_clk(flash_clk_core),
	.spimemio_flash_io0_oeb(flash_io0_oeb_core),
	.spimemio_flash_io1_oeb(flash_io1_oeb_core),
	.spimemio_flash_io2_oeb(flash_io2_oeb_core),
	.spimemio_flash_io3_oeb(flash_io3_oeb_core),
	.spimemio_flash_io0_do(flash_io0_do_core),
	.spimemio_flash_io1_do(flash_io1_do_core),
	.spimemio_flash_io2_do(flash_io2_do_core),
	.spimemio_flash_io3_do(flash_io3_do_core),
	.spimemio_flash_io0_di(flash_io0_di_core),
	.spimemio_flash_io1_di(flash_io1_di_core),
	.spimemio_flash_io2_di(flash_io2_di_core),
	.spimemio_flash_io3_di(flash_io3_di_core),

	.pad_flash_csb(flash_csb_frame),
	.pad_flash_csb_oeb(flash_csb_oeb),
	.pad_flash_clk(flash_clk_frame),
	.pad_flash_clk_oeb(flash_clk_oeb),
	.pad_flash_io0_oeb(flash_io0_oeb),
	.pad_flash_io1_oeb(flash_io1_oeb),
	.pad_flash_io0_ieb(flash_io0_ieb),
	.pad_flash_io1_ieb(flash_io1_ieb),
	.pad_flash_io0_do(flash_io0_do),
	.pad_flash_io1_do(flash_io1_do),
	.pad_flash_io0_di(flash_io0_di_buf),
	.pad_flash_io1_di(flash_io1_di_buf),








	.usr1_vcc_pwrgood(mprj_vcc_pwrgood),
	.usr2_vcc_pwrgood(mprj2_vcc_pwrgood),
	.usr1_vdd_pwrgood(mprj_vdd_pwrgood),
	.usr2_vdd_pwrgood(mprj2_vdd_pwrgood)
    );

    /* GPIO defaults (via programmed) */
    wire [((19 + 19) - (5 + 6))*13-1:0] gpio_defaults;

    /* Fixed defaults for the first 5 GPIO pins */

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h1803)
    ) gpio_defaults_block_0 (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	
	.gpio_defaults(gpio_defaults[12:0])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h1803)
    ) gpio_defaults_block_1 (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	
	.gpio_defaults(gpio_defaults[25:13])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_2 (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	
	.gpio_defaults(gpio_defaults[38:26])
    );

    // CSB is configured to be a weak pull-up
    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0801)
    ) gpio_defaults_block_3 (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	
	.gpio_defaults(gpio_defaults[51:39])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_4 (
	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
	
	.gpio_defaults(gpio_defaults[64:52])
    );

    /* Via-programmable defaults for the rest of the GPIO pins */

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_5 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[77:65])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_6 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[90:78])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_7 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[103:91])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_8 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[116:104])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_9 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[129:117])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_10 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[142:130])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_11 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[155:143])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_12 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[168:156])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_13 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[181:169])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_25 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[194:182])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_26 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[207:195])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_27 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[220:208])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_28 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[233:221])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_29 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[246:234])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_30 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[259:247])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_31 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[272:260])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_32 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[285:273])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_33 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[298:286])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_34 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[311:299])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_35 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[324:312])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_36 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[337:325])
    );

    gpio_defaults_block #(
	.GPIO_CONFIG_INIT(13'h0403)
    ) gpio_defaults_block_37 (
    	
	    .VPWR(vccd_core),
	    .VGND(vssd_core),
        
	.gpio_defaults(gpio_defaults[350:338])
    );

    // Each control block sits next to an I/O pad in the user area.
    // It gets input through a serial chain from the previous control
    // block and passes it to the next control block.  Due to the nature
    // of the shift register, bits are presented in reverse, as the first
    // bit in ends up as the last bit of the last I/O pad control block.

    // There are two types of block;  the first two and the last two
    // are configured to be full bidirectional under control of the
    // management Soc (JTAG and SDO for the first two;  flash_io2 and
    // flash_io3 for the last two).  The rest are configured to be default
    // (input).  Note that the first two and last two are the ones closest
    // to the management SoC on either side, which minimizes the wire length
    // of the extra signals those pads need.

    /* First two GPIOs (JTAG and SDO) */
    gpio_control_block gpio_control_bidir_1 [1:0] (
   	
	    .vccd(vccd_core),
	    .vssd(vssd_core),
	    .vccd1(vccd1_core),
	    .vssd1(vssd1_core),
	

	.gpio_defaults(gpio_defaults[25:0]),

    	// Management Soc-facing signals

	.resetn(gpio_resetn_1_shifted[1:0]),
	.serial_clock(gpio_clock_1_shifted[1:0]),
	.serial_load(gpio_load_1_shifted[1:0]),

	.resetn_out(gpio_resetn_1[1:0]),
	.serial_clock_out(gpio_clock_1[1:0]),
	.serial_load_out(gpio_load_1[1:0]),

    	.mgmt_gpio_in(mgmt_io_in[1:0]),
	.mgmt_gpio_out(mgmt_io_out[1:0]),
	.mgmt_gpio_oeb(mgmt_io_oeb[1:0]),

        .one(mprj_io_one[1:0]),
        .zero(mprj_io_zero[1:0]),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_1_shifted[1:0]),
    	.serial_data_out(gpio_serial_link_1[1:0]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[1:0]),
    	.user_gpio_oeb(user_io_oeb[1:0]),
    	.user_gpio_in(user_io_in[1:0]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[1:0]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[1:0]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[1:0]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[1:0]),
    	.pad_gpio_holdover(mprj_io_holdover[1:0]),
    	.pad_gpio_ana_en(mprj_io_analog_en[1:0]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[1:0]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[1:0]),
    	.pad_gpio_dm(mprj_io_dm[5:0]),
    	.pad_gpio_outenb(mprj_io_oeb[1:0]),
    	.pad_gpio_out(mprj_io_out[1:0]),
    	.pad_gpio_in(mprj_io_in[1:0])
    );

    /* Section 1 GPIOs (GPIO 0 to 18) */

    /* Section 1 GPIOs (GPIO 2 to 7) that start up under management control */

    gpio_control_block gpio_control_in_1a [5:0] (
	
            .vccd(vccd_core),
	    .vssd(vssd_core),
	    .vccd1(vccd1_core),
	    .vssd1(vssd1_core),
	

	.gpio_defaults(gpio_defaults[103:26]),

    	// Management Soc-facing signals

	.resetn(gpio_resetn_1_shifted[7:2]),
	.serial_clock(gpio_clock_1_shifted[7:2]),
	.serial_load(gpio_load_1_shifted[7:2]),

	.resetn_out(gpio_resetn_1[7:2]),
	.serial_clock_out(gpio_clock_1[7:2]),
	.serial_load_out(gpio_load_1[7:2]),

	.mgmt_gpio_in(mgmt_io_in[7:2]),
	.mgmt_gpio_out(mgmt_io_out[7:2]),
	.mgmt_gpio_oeb(mprj_io_one[7:2]),

        .one(mprj_io_one[7:2]),
        .zero(mprj_io_zero[7:2]),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_1_shifted[7:2]),
    	.serial_data_out(gpio_serial_link_1[7:2]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[7:2]),
    	.user_gpio_oeb(user_io_oeb[7:2]),
    	.user_gpio_in(user_io_in[7:2]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[7:2]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[7:2]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[7:2]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[7:2]),
    	.pad_gpio_holdover(mprj_io_holdover[7:2]),
    	.pad_gpio_ana_en(mprj_io_analog_en[7:2]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[7:2]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[7:2]),
    	.pad_gpio_dm(mprj_io_dm[23:6]),
    	.pad_gpio_outenb(mprj_io_oeb[7:2]),
    	.pad_gpio_out(mprj_io_out[7:2]),
    	.pad_gpio_in(mprj_io_in[7:2])
    );

    /* Section 1 GPIOs (GPIO 8 to 18) */
    gpio_control_block gpio_control_in_1 [19-5-9:0] (
	
            .vccd(vccd_core),
	    .vssd(vssd_core),
	    .vccd1(vccd1_core),
	    .vssd1(vssd1_core),
	

	.gpio_defaults(gpio_defaults[((19-5)*13-1):104]),

    	// Management Soc-facing signals

	.resetn(gpio_resetn_1_shifted[(19-5-1):8]),
	.serial_clock(gpio_clock_1_shifted[(19-5-1):8]),
	.serial_load(gpio_load_1_shifted[(19-5-1):8]),

	.resetn_out(gpio_resetn_1[(19-5-1):8]),
	.serial_clock_out(gpio_clock_1[(19-5-1):8]),
	.serial_load_out(gpio_load_1[(19-5-1):8]),

	.mgmt_gpio_in(mgmt_io_in[(19 - 5 - 1):8]),
	.mgmt_gpio_out(mgmt_io_out[(19 - 5 - 1):8]),
	.mgmt_gpio_oeb(mprj_io_one[(19-5-1):8]),
  
        .one(mprj_io_one[(19-5-1):8]),
        .zero(),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_1_shifted[(19-5-1):8]),
    	.serial_data_out(gpio_serial_link_1[(19-5-1):8]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[(19-5-1):8]),
    	.user_gpio_oeb(user_io_oeb[(19-5-1):8]),
    	.user_gpio_in(user_io_in[(19-5-1):8]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[(19-5-1):8]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[(19-5-1):8]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[(19-5-1):8]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[(19-5-1):8]),
    	.pad_gpio_holdover(mprj_io_holdover[(19-5-1):8]),
    	.pad_gpio_ana_en(mprj_io_analog_en[(19-5-1):8]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[(19-5-1):8]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[(19-5-1):8]),
    	.pad_gpio_dm(mprj_io_dm[(19-5)*3-1:24]),
    	.pad_gpio_outenb(mprj_io_oeb[(19-5-1):8]),
    	.pad_gpio_out(mprj_io_out[(19-5-1):8]),
    	.pad_gpio_in(mprj_io_in[(19-5-1):8])
    );

    /* Last three GPIOs (spi_sdo, flash_io2 and flash_io3) */

    gpio_control_block gpio_control_bidir_2 [2:0] (
    	
	    .vccd(vccd_core),
	    .vssd(vssd_core),
	    .vccd1(vccd1_core),
	    .vssd1(vssd1_core),
        

	.gpio_defaults(gpio_defaults[(((19 + 19)-(5 + 6))*13-1):(((19 + 19)-(5 + 6))*13-39)]),

    	// Management Soc-facing signals

	.resetn(gpio_resetn_2_shifted[(19-6-1):(19-6-3)]),
	.serial_clock(gpio_clock_2_shifted[(19-6-1):(19-6-3)]),
	.serial_load(gpio_load_2_shifted[(19-6-1):(19-6-3)]),

	.resetn_out(gpio_resetn_2[(19-6-1):(19-6-3)]),
	.serial_clock_out(gpio_clock_2[(19-6-1):(19-6-3)]),
	.serial_load_out(gpio_load_2[(19-6-1):(19-6-3)]),

	.mgmt_gpio_in(mgmt_io_in[(((19 + 19) - 1)):(((19 + 19) - 1)-2)]),
	.mgmt_gpio_out(mgmt_io_out[(((19 + 19) - 1)):(((19 + 19) - 1)-2)]),
	.mgmt_gpio_oeb(mgmt_io_oeb[(((19 + 19) - 1)):(((19 + 19) - 1)-2)]),

        .one(mprj_io_one[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
        .zero(),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_2_shifted[(19-6-1):(19-6-3)]),
    	.serial_data_out(gpio_serial_link_2[(19-6-1):(19-6-3)]),

    	// User-facing signals
    	.user_gpio_out(user_io_out[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.user_gpio_oeb(user_io_oeb[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.user_gpio_in(user_io_in[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_holdover(mprj_io_holdover[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_ana_en(mprj_io_analog_en[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_dm(mprj_io_dm[(((19 + 19) - (5 + 6))*3-1):(((19 + 19) - (5 + 6))*3-9)]),
    	.pad_gpio_outenb(mprj_io_oeb[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_out(mprj_io_out[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)]),
    	.pad_gpio_in(mprj_io_in[(((19 + 19) - (5 + 6))-1):(((19 + 19) - (5 + 6))-3)])
    );

    /* Section 2 GPIOs (GPIO 19 to 37) */

    gpio_control_block gpio_control_in_2 [19-6-4:0] (
	
            .vccd(vccd_core),
	    .vssd(vssd_core),
	    .vccd1(vccd1_core),
	    .vssd1(vssd1_core),
	

 	.gpio_defaults(gpio_defaults[(((19 + 19)-(5 + 6)-3)*13-1):((19-5)*13)]),

    	// Management Soc-facing signals

	.resetn(gpio_resetn_2_shifted[(19-6-4):0]),
	.serial_clock(gpio_clock_2_shifted[(19-6-4):0]),
	.serial_load(gpio_load_2_shifted[(19-6-4):0]),

	.resetn_out(gpio_resetn_2[(19-6-4):0]),
	.serial_clock_out(gpio_clock_2[(19-6-4):0]),
	.serial_load_out(gpio_load_2[(19-6-4):0]),

 	.mgmt_gpio_in(mgmt_io_in[(((19 + 19) - 1)-3):(19 + 6)]),
 	.mgmt_gpio_out(mgmt_io_out[(((19 + 19) - 1)-3):(19 + 6)]),
	.mgmt_gpio_oeb(mprj_io_one[(((19 + 19) - (5 + 6))-4):(19-5)]),
	.one(mprj_io_one[(((19 + 19) - (5 + 6))-4):(19-5)]),
        .zero(),

    	// Serial data chain for pad configuration
    	.serial_data_in(gpio_serial_link_2_shifted[(19-6-4):0]),
    	.serial_data_out(gpio_serial_link_2[(19-6-4):0]),

    	// User-facing signals
   	.user_gpio_out(user_io_out[(((19 + 19) - (5 + 6))-4):(19-5)]),
   	.user_gpio_oeb(user_io_oeb[(((19 + 19) - (5 + 6))-4):(19-5)]),
  	.user_gpio_in(user_io_in[(((19 + 19) - (5 + 6))-4):(19-5)]),

    	// Pad-facing signals (Pad GPIOv2)
    	.pad_gpio_inenb(mprj_io_inp_dis[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_ib_mode_sel(mprj_io_ib_mode_sel[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_vtrip_sel(mprj_io_vtrip_sel[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_slow_sel(mprj_io_slow_sel[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_holdover(mprj_io_holdover[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_ana_en(mprj_io_analog_en[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_ana_sel(mprj_io_analog_sel[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_ana_pol(mprj_io_analog_pol[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_dm(mprj_io_dm[((((19 + 19) - (5 + 6)))*3-10):((19-5)*3)]),
    	.pad_gpio_outenb(mprj_io_oeb[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_out(mprj_io_out[(((19 + 19) - (5 + 6))-4):(19-5)]),
    	.pad_gpio_in(mprj_io_in[(((19 + 19) - (5 + 6))-4):(19-5)])
    );

    user_id_programming #(
	.USER_PROJECT_ID(USER_PROJECT_ID)
    ) user_id_value (
	
		.VPWR(vccd_core),
		.VGND(vssd_core),
	
	.mask_rev(mask_rev)
    );

    // Power-on-reset circuit
    simple_por por (
	
		.vdd3v3(vddio_core),
		.vdd1v8(vccd_core),
		.vss3v3(vssio_core),
		.vss1v8(vssd_core),
	
		.porb_h(porb_h),
		.porb_l(porb_l),
		.por_l(por_l)
    );

    // XRES (chip input pin reset) reset level converter
    xres_buf rstb_level (
	
		.VPWR(vddio_core),
		.LVPWR(vccd_core),
		.LVGND(vssd_core),
		.VGND(vssio_core),
	
		.A(rstb_h),
		.X(rstb_l)
    );

    /* Spare logic for metal mask fixes */
    // `define NUM_SPARE_BLOCKS (`MPRJ_DIG_PADS+4)
    

    wire [(27*4)-1:0] spare_xz_nc;
    wire [(4*4)-1:0] spare_xi_nc;
    wire [(1*4)-1:0] spare_xib_nc;
    wire [(2*4)-1:0] spare_xna_nc;
    wire [(2*4)-1:0] spare_xno_nc;
    wire [(2*4)-1:0] spare_xmx_nc;
    wire [(2*4)-1:0] spare_xfq_nc;
    wire [(2*4)-1:0] spare_xfqn_nc;

    // Four spare logic blocks above the processor and one per GPIO
    // control block.
    spare_logic_block spare_logic [4-1:0] (
	
		.vccd(vccd_core),
		.vssd(vssd_core),
	
		.spare_xz(spare_xz_nc),
		.spare_xi(spare_xi_nc),
		.spare_xib(spare_xib_nc),
		.spare_xna(spare_xna_nc),
		.spare_xno(spare_xno_nc),
		.spare_xmx(spare_xmx_nc),
		.spare_xfq(spare_xfq_nc),
		.spare_xfqn(spare_xfqn_nc)
    );

    









endmodule
// `default_nettype wire
module empty_macro ();
endmodule
module manual_power_connections ();
endmodule
module copyright_block ();
endmodule
module caravel_logo ();
endmodule
module caravel_motto ();
endmodule
module open_source ();
endmodule
module user_id_textblock ();
endmodule
module gpio_defaults_block_0403 (VGND,
    VPWR,
    gpio_defaults);
 input VGND;
 input VPWR;
 output [12:0] gpio_defaults;

 wire \gpio_defaults_low[0] ;
 wire \gpio_defaults_high[10] ;
 wire \gpio_defaults_low[11] ;
 wire \gpio_defaults_low[12] ;
 wire \gpio_defaults_high[1] ;
 wire \gpio_defaults_low[2] ;
 wire \gpio_defaults_low[3] ;
 wire \gpio_defaults_low[4] ;
 wire \gpio_defaults_low[5] ;
 wire \gpio_defaults_low[6] ;
 wire \gpio_defaults_low[7] ;
 wire \gpio_defaults_low[8] ;
 wire \gpio_defaults_low[9] ;
 wire \gpio_defaults_high[0] ;
 wire \gpio_defaults_high[11] ;
 wire \gpio_defaults_high[12] ;
 wire \gpio_defaults_high[2] ;
 wire \gpio_defaults_high[3] ;
 wire \gpio_defaults_high[4] ;
 wire \gpio_defaults_high[5] ;
 wire \gpio_defaults_high[6] ;
 wire \gpio_defaults_high[7] ;
 wire \gpio_defaults_high[8] ;
 wire \gpio_defaults_high[9] ;
 wire \gpio_defaults_low[10] ;
 wire \gpio_defaults_low[1] ;

 sky130_fd_sc_hd__fill_1 FILLER_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[0]  (.HI(\gpio_defaults_high[0] ),
    .LO(\gpio_defaults_low[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[10]  (.HI(\gpio_defaults_high[10] ),
    .LO(\gpio_defaults_low[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[11]  (.HI(\gpio_defaults_high[11] ),
    .LO(\gpio_defaults_low[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[12]  (.HI(\gpio_defaults_high[12] ),
    .LO(\gpio_defaults_low[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[1]  (.HI(\gpio_defaults_high[1] ),
    .LO(\gpio_defaults_low[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[2]  (.HI(\gpio_defaults_high[2] ),
    .LO(\gpio_defaults_low[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[3]  (.HI(\gpio_defaults_high[3] ),
    .LO(\gpio_defaults_low[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[4]  (.HI(\gpio_defaults_high[4] ),
    .LO(\gpio_defaults_low[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[5]  (.HI(\gpio_defaults_high[5] ),
    .LO(\gpio_defaults_low[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[6]  (.HI(\gpio_defaults_high[6] ),
    .LO(\gpio_defaults_low[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[7]  (.HI(\gpio_defaults_high[7] ),
    .LO(\gpio_defaults_low[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[8]  (.HI(\gpio_defaults_high[8] ),
    .LO(\gpio_defaults_low[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[9]  (.HI(\gpio_defaults_high[9] ),
    .LO(\gpio_defaults_low[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign gpio_defaults[0] = \gpio_defaults_high[0] ;
 assign gpio_defaults[1] = \gpio_defaults_high[1] ;
 assign gpio_defaults[2] = \gpio_defaults_low[2] ;
 assign gpio_defaults[3] = \gpio_defaults_low[3] ;
 assign gpio_defaults[4] = \gpio_defaults_low[4] ;
 assign gpio_defaults[5] = \gpio_defaults_low[5] ;
 assign gpio_defaults[6] = \gpio_defaults_low[6] ;
 assign gpio_defaults[7] = \gpio_defaults_low[7] ;
 assign gpio_defaults[8] = \gpio_defaults_low[8] ;
 assign gpio_defaults[9] = \gpio_defaults_low[9] ;
 assign gpio_defaults[10] = \gpio_defaults_high[10] ;
 assign gpio_defaults[11] = \gpio_defaults_low[11] ;
 assign gpio_defaults[12] = \gpio_defaults_low[12] ;
endmodule
module gpio_defaults_block_1803 (VGND,
    VPWR,
    gpio_defaults);
 input VGND;
 input VPWR;
 output [12:0] gpio_defaults;

 wire \gpio_defaults_low[0] ;
 wire \gpio_defaults_high[10] ;
 wire \gpio_defaults_low[11] ;
 wire \gpio_defaults_low[12] ;
 wire \gpio_defaults_high[1] ;
 wire \gpio_defaults_low[2] ;
 wire \gpio_defaults_low[3] ;
 wire \gpio_defaults_low[4] ;
 wire \gpio_defaults_low[5] ;
 wire \gpio_defaults_low[6] ;
 wire \gpio_defaults_low[7] ;
 wire \gpio_defaults_low[8] ;
 wire \gpio_defaults_low[9] ;
 wire \gpio_defaults_high[0] ;
 wire \gpio_defaults_high[11] ;
 wire \gpio_defaults_high[12] ;
 wire \gpio_defaults_high[2] ;
 wire \gpio_defaults_high[3] ;
 wire \gpio_defaults_high[4] ;
 wire \gpio_defaults_high[5] ;
 wire \gpio_defaults_high[6] ;
 wire \gpio_defaults_high[7] ;
 wire \gpio_defaults_high[8] ;
 wire \gpio_defaults_high[9] ;
 wire \gpio_defaults_low[10] ;
 wire \gpio_defaults_low[1] ;

 sky130_fd_sc_hd__fill_1 FILLER_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[0]  (.HI(\gpio_defaults_high[0] ),
    .LO(\gpio_defaults_low[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[10]  (.HI(\gpio_defaults_high[10] ),
    .LO(\gpio_defaults_low[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[11]  (.HI(\gpio_defaults_high[11] ),
    .LO(\gpio_defaults_low[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[12]  (.HI(\gpio_defaults_high[12] ),
    .LO(\gpio_defaults_low[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[1]  (.HI(\gpio_defaults_high[1] ),
    .LO(\gpio_defaults_low[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[2]  (.HI(\gpio_defaults_high[2] ),
    .LO(\gpio_defaults_low[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[3]  (.HI(\gpio_defaults_high[3] ),
    .LO(\gpio_defaults_low[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[4]  (.HI(\gpio_defaults_high[4] ),
    .LO(\gpio_defaults_low[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[5]  (.HI(\gpio_defaults_high[5] ),
    .LO(\gpio_defaults_low[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[6]  (.HI(\gpio_defaults_high[6] ),
    .LO(\gpio_defaults_low[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[7]  (.HI(\gpio_defaults_high[7] ),
    .LO(\gpio_defaults_low[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[8]  (.HI(\gpio_defaults_high[8] ),
    .LO(\gpio_defaults_low[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[9]  (.HI(\gpio_defaults_high[9] ),
    .LO(\gpio_defaults_low[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign gpio_defaults[0] = \gpio_defaults_high[0] ;
 assign gpio_defaults[1] = \gpio_defaults_high[1] ;
 assign gpio_defaults[2] = \gpio_defaults_low[2] ;
 assign gpio_defaults[3] = \gpio_defaults_low[3] ;
 assign gpio_defaults[4] = \gpio_defaults_low[4] ;
 assign gpio_defaults[5] = \gpio_defaults_low[5] ;
 assign gpio_defaults[6] = \gpio_defaults_low[6] ;
 assign gpio_defaults[7] = \gpio_defaults_low[7] ;
 assign gpio_defaults[8] = \gpio_defaults_low[8] ;
 assign gpio_defaults[9] = \gpio_defaults_low[9] ;
 assign gpio_defaults[10] = \gpio_defaults_low[10] ;
 assign gpio_defaults[11] = \gpio_defaults_high[11] ;
 assign gpio_defaults[12] = \gpio_defaults_high[12] ;
endmodule
module gpio_defaults_block_0801 (VGND,
    VPWR,
    gpio_defaults);
 input VGND;
 input VPWR;
 output [12:0] gpio_defaults;

 wire \gpio_defaults_low[0] ;
 wire \gpio_defaults_high[10] ;
 wire \gpio_defaults_low[11] ;
 wire \gpio_defaults_low[12] ;
 wire \gpio_defaults_high[1] ;
 wire \gpio_defaults_low[2] ;
 wire \gpio_defaults_low[3] ;
 wire \gpio_defaults_low[4] ;
 wire \gpio_defaults_low[5] ;
 wire \gpio_defaults_low[6] ;
 wire \gpio_defaults_low[7] ;
 wire \gpio_defaults_low[8] ;
 wire \gpio_defaults_low[9] ;
 wire \gpio_defaults_high[0] ;
 wire \gpio_defaults_high[11] ;
 wire \gpio_defaults_high[12] ;
 wire \gpio_defaults_high[2] ;
 wire \gpio_defaults_high[3] ;
 wire \gpio_defaults_high[4] ;
 wire \gpio_defaults_high[5] ;
 wire \gpio_defaults_high[6] ;
 wire \gpio_defaults_high[7] ;
 wire \gpio_defaults_high[8] ;
 wire \gpio_defaults_high[9] ;
 wire \gpio_defaults_low[10] ;
 wire \gpio_defaults_low[1] ;

 sky130_fd_sc_hd__fill_1 FILLER_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[0]  (.HI(\gpio_defaults_high[0] ),
    .LO(\gpio_defaults_low[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[10]  (.HI(\gpio_defaults_high[10] ),
    .LO(\gpio_defaults_low[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[11]  (.HI(\gpio_defaults_high[11] ),
    .LO(\gpio_defaults_low[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[12]  (.HI(\gpio_defaults_high[12] ),
    .LO(\gpio_defaults_low[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[1]  (.HI(\gpio_defaults_high[1] ),
    .LO(\gpio_defaults_low[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[2]  (.HI(\gpio_defaults_high[2] ),
    .LO(\gpio_defaults_low[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[3]  (.HI(\gpio_defaults_high[3] ),
    .LO(\gpio_defaults_low[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[4]  (.HI(\gpio_defaults_high[4] ),
    .LO(\gpio_defaults_low[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[5]  (.HI(\gpio_defaults_high[5] ),
    .LO(\gpio_defaults_low[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[6]  (.HI(\gpio_defaults_high[6] ),
    .LO(\gpio_defaults_low[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[7]  (.HI(\gpio_defaults_high[7] ),
    .LO(\gpio_defaults_low[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[8]  (.HI(\gpio_defaults_high[8] ),
    .LO(\gpio_defaults_low[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[9]  (.HI(\gpio_defaults_high[9] ),
    .LO(\gpio_defaults_low[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign gpio_defaults[0] = \gpio_defaults_high[0] ;
 assign gpio_defaults[1] = \gpio_defaults_low[1] ;
 assign gpio_defaults[2] = \gpio_defaults_low[2] ;
 assign gpio_defaults[3] = \gpio_defaults_low[3] ;
 assign gpio_defaults[4] = \gpio_defaults_low[4] ;
 assign gpio_defaults[5] = \gpio_defaults_low[5] ;
 assign gpio_defaults[6] = \gpio_defaults_low[6] ;
 assign gpio_defaults[7] = \gpio_defaults_low[7] ;
 assign gpio_defaults[8] = \gpio_defaults_low[8] ;
 assign gpio_defaults[9] = \gpio_defaults_low[9] ;
 assign gpio_defaults[10] = \gpio_defaults_low[10] ;
 assign gpio_defaults[11] = \gpio_defaults_high[11] ;
 assign gpio_defaults[12] = \gpio_defaults_low[12] ;
endmodule
/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_gpio_ovtv2: General Purpose I/0.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_gpio_ovtv2 ( IN, IN_H, TIE_HI_ESD, TIE_LO_ESD, AMUXBUS_A,
                                      AMUXBUS_B, PAD, PAD_A_ESD_0_H, PAD_A_ESD_1_H, PAD_A_NOESD_H,
                                      VCCD, VCCHIB,VDDA, VDDIO, VDDIO_Q, VSSA, VSSD, VSSIO, VSSIO_Q, VSWITCH,
                                      ANALOG_EN, ANALOG_POL, ANALOG_SEL, DM, ENABLE_H, ENABLE_INP_H, ENABLE_VDDA_H, ENABLE_VDDIO, ENABLE_VSWITCH_H, HLD_H_N,
                                      HLD_OVR, IB_MODE_SEL, INP_DIS, OE_N, OUT, SLOW, SLEW_CTL, VTRIP_SEL, HYS_TRIM, VINREF );
input OUT;
input OE_N;
input HLD_H_N;
input ENABLE_H;
input ENABLE_INP_H;
input ENABLE_VDDA_H;
input ENABLE_VDDIO;
input ENABLE_VSWITCH_H;
input INP_DIS;
input VTRIP_SEL;
input HYS_TRIM;
input SLOW;
input [1:0] SLEW_CTL;
input HLD_OVR;
input ANALOG_EN;
input ANALOG_SEL;
input ANALOG_POL;
input [2:0] DM;
input [1:0] IB_MODE_SEL;
input VINREF;
inout VDDIO;
inout VDDIO_Q;
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;
inout PAD;
inout PAD_A_NOESD_H,PAD_A_ESD_0_H,PAD_A_ESD_1_H;
inout AMUXBUS_A;
inout AMUXBUS_B;
output IN;
output IN_H;
output TIE_HI_ESD, TIE_LO_ESD;
wire hld_h_n_del;
wire hld_h_n_buf;
reg [2:0] dm_final;
reg [1:0] slew_ctl_final;
reg slow_final, vtrip_sel_final, inp_dis_final, out_final, oe_n_final, hld_ovr_final, hys_trim_final, analog_en_final,analog_en_vdda, analog_en_vswitch,analog_en_vddio_q;
reg [1:0] ib_mode_sel_final;
wire [2:0] dm_del;
wire [1:0] slew_ctl_del;
wire [1:0] ib_mode_sel_del;
wire slow_del, vtrip_sel_del, inp_dis_del, out_del, oe_n_del, hld_ovr_del, hys_trim_del;
wire [2:0] dm_buf;
wire [1:0] slew_ctl_buf;
wire [1:0] ib_mode_sel_buf;
wire slow_buf, vtrip_sel_buf, inp_dis_buf, out_buf, oe_n_buf, hld_ovr_buf, hys_trim_buf;
reg notifier_dm, notifier_slow, notifier_oe_n, notifier_out, notifier_vtrip_sel, notifier_hld_ovr, notifier_inp_dis;
reg notifier_slew_ctl, notifier_ib_mode_sel, notifier_hys_trim;
reg notifier_enable_h, notifier, dummy_notifier1;
assign hld_h_n_buf 	= HLD_H_N;
assign hld_ovr_buf 	= HLD_OVR;
assign dm_buf 		= DM;
assign inp_dis_buf 	= INP_DIS;
assign vtrip_sel_buf 	= VTRIP_SEL;
assign slow_buf 	= SLOW;
assign oe_n_buf 	= OE_N;
assign out_buf 		= OUT;
assign ib_mode_sel_buf 	= IB_MODE_SEL;
assign slew_ctl_buf	= SLEW_CTL;
assign hys_trim_buf 	= HYS_TRIM;
wire  pwr_good_amux	         = ((hld_h_n_buf===0 || ENABLE_H===0) ? 1:(VCCD===1))  && (VSSD===0) && (VSSA===0) && (VSSIO_Q===0);
wire  pwr_good_output_driver     = (VDDIO===1)   && (VDDIO_Q===1)&& (VSSIO===0)   && (VSSD===0)  && (VSSA===0) ;
wire  pwr_good_hold_ovr_mode     = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0)    && (VCCHIB===1);
wire  pwr_good_active_mode       = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0)    && (VCCD===1);
wire  pwr_good_hold_mode         = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0);
wire  pwr_good_active_mode_vdda  = (VDDA===1)  && (VSSD===0)   && (VCCD===1);
wire  pwr_good_hold_mode_vdda    = (VDDA===1)    && (VSSD===0);
wire  pwr_good_inpbuff_hv        = (VDDIO_Q===1) && (inp_dis_final===0 && dm_final!==3'b000 && ib_mode_sel_final===2'b01 ? VCCHIB===1 : 1) && (VSSD===0);
wire  pwr_good_inpbuff_lv        = (VDDIO_Q===1) && (VSSD===0)   && (VCCHIB===1);
wire  pwr_good_analog_en_vdda    = (VDDA===1)  && (VSSD===0) && (VSSA===0) ;
wire  pwr_good_analog_en_vddio_q = (VDDIO_Q ===1)  && (VSSD===0) && (VSSA===0) ;
wire  pwr_good_analog_en_vswitch = (VSWITCH ===1)  && (VSSD===0) && (VSSA===0) ;
wire  pwr_good_amux_vccd   	 = ((hld_h_n_buf===0 || ENABLE_H===0) ? 1:(VCCD===1));
parameter MAX_WARNING_COUNT = 100;
wire pad_tristate = oe_n_final === 1 || dm_final === 3'b000 || dm_final === 3'b001;
wire x_on_pad  =  !pwr_good_output_driver
     || (dm_final !== 3'b000 	&& dm_final !== 3'b001 		&& oe_n_final===1'bx)
     || (^dm_final[2:0] === 1'bx 	&& oe_n_final===1'b0)
     || (slow_final===1'bx 	&& dm_final !== 3'b000		&& dm_final !== 3'b001 && oe_n_final===1'b0)
     || (slow_final===1'b1 	&& ^slew_ctl_final[1:0] ===1'bx 	&& dm_final === 3'b100 && oe_n_final===1'b0);




parameter SLOW_1_DELAY= 0;
parameter SLOW_0_DELAY= 0;







parameter SLEW_00_DELAY= 0 ;
parameter SLEW_01_DELAY= 0;
parameter SLEW_10_DELAY= 0;
parameter SLEW_11_DELAY= 0;

integer slow_1_delay,slow_0_delay,slow_delay,slew_00_delay,slew_01_delay,slew_10_delay,slew_11_delay;
initial slow_1_delay = SLOW_1_DELAY;
initial slow_0_delay = SLOW_0_DELAY;
initial slew_00_delay = SLEW_00_DELAY;
initial slew_01_delay = SLEW_01_DELAY;
initial slew_10_delay = SLEW_10_DELAY;
initial slew_11_delay = SLEW_11_DELAY;
always @(*)
begin
    if (SLOW===1)
    begin
        if (DM[2]===1 && DM[1]===0 && DM[0]===0)
        begin










            slow_delay = slow_1_delay;

        end
        else
            slow_delay = slow_1_delay;
    end
    else
        slow_delay = slow_0_delay;
end
bufif1 (pull1, strong0) #slow_delay dm2 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b010));
bufif1 (strong1, pull0) #slow_delay dm3 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b011));
bufif1 (highz1, strong0) #slow_delay dm4 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b100));
bufif1 (strong1, highz0) #slow_delay dm5 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b101));
bufif1 (strong1, strong0) #slow_delay dm6 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b110));
bufif1 (pull1, pull0)  #slow_delay dm7 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b111));
tran pad_esd_1 (PAD,PAD_A_NOESD_H);
tran pad_esd_2 (PAD,PAD_A_ESD_0_H);
tran pad_esd_3 (PAD,PAD_A_ESD_1_H);
wire x_on_in_hv  =  (ENABLE_H===0  && ^ENABLE_INP_H===1'bx)
     || (inp_dis_final===1'bx  && ^dm_final[2:0]!==1'bx && dm_final !== 3'b000)
     || (^ENABLE_H===1'bx)
     || (inp_dis_final===0 	       		&& ^dm_final[2:0] === 1'bx)
     || (^ib_mode_sel_final===1'bx  	&& inp_dis_final===0  		&& dm_final !== 3'b000)
     || (vtrip_sel_final===1'bx    		&& inp_dis_final===0        	&& dm_final !== 3'b000		&& ib_mode_sel_final===2'b00)
     || (^ENABLE_VDDIO===1'bx    		&& inp_dis_final===0        	&& dm_final !== 3'b000		&& ib_mode_sel_final===2'b01)
     || (ib_mode_sel_final[1]===1'b1	&& VINREF !== 1'b1    		&& inp_dis_final===0      	&& dm_final !== 3'b000)
     || (ib_mode_sel_final[1]===1'b1	&& hys_trim_final===1'bx	&& inp_dis_final===0      	&& dm_final !== 3'b000);
wire x_on_in_lv  =  (ENABLE_H===0  && ^ENABLE_VDDIO===1'bx)
     || (ENABLE_H===0  && ^ENABLE_INP_H===1'bx)
     || (inp_dis_final===1'bx  && ^dm_final[2:0]!==1'bx && dm_final !== 3'b000)
     || (^ENABLE_H===1'bx)
     || (inp_dis_final===0 	       		&& ^dm_final[2:0] === 1'bx)
     || (^ib_mode_sel_final===1'bx  	&& inp_dis_final===0  		&& dm_final !== 3'b000)
     || (vtrip_sel_final===1'bx    		&& inp_dis_final===0        	&& dm_final !== 3'b000		&& ib_mode_sel_final===2'b00)
     || (^ENABLE_VDDIO===1'bx    		&& inp_dis_final===0        	&& dm_final !== 3'b000	)
     || (ib_mode_sel_final[1]===1'b1	&& VINREF !== 1'b1    		&& inp_dis_final===0      	&& dm_final !== 3'b000)
     || (ib_mode_sel_final[1]===1'b1	&& hys_trim_final===1'bx	&& inp_dis_final===0      	&& dm_final !== 3'b000);
wire disable_inp_buff = ENABLE_H===1 ? (dm_final===3'b000 || inp_dis_final===1) : ENABLE_INP_H===0;
assign IN_H = (x_on_in_hv===1 || pwr_good_inpbuff_hv===0) ? 1'bx : (disable_inp_buff===1 ? 0 : (^PAD===1'bx ? 1'bx : PAD));
wire disable_inp_buff_lv = ENABLE_H===1 ? (dm_final===3'b000 || inp_dis_final===1) : ENABLE_VDDIO===0;
assign IN   = (x_on_in_lv ===1 || pwr_good_inpbuff_lv===0) ? 1'bx : (disable_inp_buff_lv===1 ? 0 : (^PAD===1'bx ? 1'bx : PAD));
assign TIE_HI_ESD = VDDIO===1'b1 ? 1'b1 : 1'bx;
assign TIE_LO_ESD = VSSIO===1'b0 ? 1'b0 : 1'bx;
wire functional_mode_amux = (pwr_good_analog_en_vdda ===1 && pwr_good_analog_en_vddio_q ===1 && pwr_good_analog_en_vswitch ===1 );
wire x_on_analog_en_vdda = (pwr_good_analog_en_vdda !==1
                            || (functional_mode_amux ==1 && (ENABLE_H !==0 && ^hld_h_n_buf === 1'bx) || (hld_h_n_buf!== 0 && ^ENABLE_H=== 1'bx) || pwr_good_amux_vccd !==1 )
                            || (functional_mode_amux ==1 && (hld_h_n_buf ===1 && ENABLE_H===1 && ^ANALOG_EN === 1'bx && ENABLE_VDDA_H ===1 && ENABLE_VSWITCH_H===1 ) || (hld_h_n_buf ===1 && ENABLE_H===1 && ANALOG_EN ===0 && ^ENABLE_VDDA_H ===1'bx) ));
wire zero_on_analog_en_vdda = ( (pwr_good_analog_en_vdda ===1 && ENABLE_VDDA_H ===0)
                                || (pwr_good_analog_en_vdda ===1 && pwr_good_analog_en_vddio_q ===1 && hld_h_n_buf===0)
                                || (pwr_good_analog_en_vdda ===1 && pwr_good_analog_en_vddio_q ===1 && ENABLE_H===0)
                                ||  (pwr_good_analog_en_vdda ===1 && pwr_good_analog_en_vddio_q ===1 && pwr_good_amux_vccd && ANALOG_EN===0) );
wire x_on_analog_en_vddio_q =  ( pwr_good_analog_en_vddio_q !==1
                                 || (functional_mode_amux ==1 && (ENABLE_H !==0 && ^hld_h_n_buf === 1'bx) || (hld_h_n_buf!== 0 && ^ENABLE_H=== 1'bx) || pwr_good_amux_vccd !==1 )
                                 || (functional_mode_amux ==1 && (hld_h_n_buf ===1 && ENABLE_H===1 && ^ANALOG_EN === 1'bx && ENABLE_VDDA_H ===1 && ENABLE_VSWITCH_H===1 ) ));
wire zero_on_analog_en_vddio_q =  ( (pwr_good_analog_en_vddio_q ===1 && hld_h_n_buf===0)
                                    || (pwr_good_analog_en_vddio_q ===1 && ENABLE_H===0)
                                    ||  (pwr_good_analog_en_vddio_q ===1 && pwr_good_amux_vccd && ANALOG_EN===0) );
wire x_on_analog_en_vswitch = (pwr_good_analog_en_vswitch !==1
                               || (functional_mode_amux ==1 && (ENABLE_H !==0 && ^hld_h_n_buf === 1'bx) || (hld_h_n_buf!== 0 && ^ENABLE_H=== 1'bx) || pwr_good_amux_vccd !==1 )
                               || (functional_mode_amux ==1 && (hld_h_n_buf ===1 && ENABLE_H===1 && ^ANALOG_EN === 1'bx && ENABLE_VDDA_H ===1 && ENABLE_VSWITCH_H===1 ) || (hld_h_n_buf ===1 && ENABLE_H===1 && ANALOG_EN ===0 && ^ENABLE_VSWITCH_H ===1'bx) ));
wire  zero_on_analog_en_vswitch =   ( (pwr_good_analog_en_vswitch ===1 && ENABLE_VSWITCH_H ===0)
                                      || (pwr_good_analog_en_vswitch ===1 && pwr_good_analog_en_vddio_q ===1 && hld_h_n_buf===0)
                                      || (pwr_good_analog_en_vswitch ===1 && pwr_good_analog_en_vddio_q ===1 && ENABLE_H===0)
                                      ||  (pwr_good_analog_en_vswitch ===1 && pwr_good_analog_en_vddio_q ===1 && pwr_good_amux_vccd && ANALOG_EN===0) );
always @(*)
begin : LATCH_dm
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        dm_final 	<= 3'bxxx;
    end
    else if (ENABLE_H===0)
    begin
        dm_final 	<= 3'b000;
    end
    else if (hld_h_n_buf===1)
    begin
        dm_final 	<= (^dm_buf[2:0]	=== 1'bx	|| !pwr_good_active_mode) ? 3'bxxx : dm_buf;
    end
end
always @(notifier_enable_h or notifier_dm)
begin
    disable LATCH_dm; dm_final <= 3'bxxx;
end
always @(*)
begin : LATCH_inp_dis
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        inp_dis_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        inp_dis_final 	<= 1'b1;
    end
    else if (hld_h_n_buf===1)
    begin
        inp_dis_final 	<= (^inp_dis_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : inp_dis_buf;
    end
end
always @(notifier_enable_h or notifier_inp_dis)
begin
    disable LATCH_inp_dis; inp_dis_final <= 1'bx;
end
always @(*)
begin : LATCH_ib_mode_sel
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        ib_mode_sel_final 	<= 2'bxx;
    end
    else if (ENABLE_H===0)
    begin
        ib_mode_sel_final 	<= 2'b00;
    end
    else if (hld_h_n_buf===1)
    begin
        ib_mode_sel_final 	<= (^ib_mode_sel_buf[1:0]	=== 1'bx	|| !pwr_good_active_mode) ? 2'bxx : ib_mode_sel_buf;
    end
end
always @(notifier_enable_h or notifier_ib_mode_sel)
begin
    disable LATCH_ib_mode_sel; ib_mode_sel_final <= 2'bxx;
end
always @(*)
begin : LATCH_slew_ctl_final
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        slew_ctl_final 	<= 2'bxx;
    end
    else if (ENABLE_H===0)
    begin
        slew_ctl_final 	<= 2'b00;
    end
    else if (hld_h_n_buf===1)
    begin
        slew_ctl_final 	<= (^slew_ctl_buf[1:0] === 1'bx || !pwr_good_active_mode) ? 2'bxx : slew_ctl_buf;
    end
end
always @(notifier_enable_h or notifier_slew_ctl)
begin
    disable LATCH_slew_ctl_final; slew_ctl_final <= 2'bxx;
end
always @(*)
begin : LATCH_vtrip_sel
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        vtrip_sel_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        vtrip_sel_final 	<= 1'b0;
    end
    else if (hld_h_n_buf===1)
    begin
        vtrip_sel_final 	<= (^vtrip_sel_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : vtrip_sel_buf;
    end
end
always @(notifier_enable_h or notifier_vtrip_sel)
begin
    disable LATCH_vtrip_sel; vtrip_sel_final <= 1'bx;
end
always @(*)
begin : LATCH_hys_trim
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        hys_trim_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        hys_trim_final 	<= 1'b0;
    end
    else if (hld_h_n_buf===1)
    begin
        hys_trim_final 	<= (^hys_trim_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : hys_trim_buf;
    end
end
always @(notifier_enable_h or notifier_hys_trim)
begin
    disable LATCH_hys_trim; hys_trim_final <= 1'bx;
end
always @(*)
begin : LATCH_slow
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        slow_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        slow_final 	<= 1'b0;
    end
    else if (hld_h_n_buf===1)
    begin
        slow_final 	<= (^slow_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : slow_buf;
    end
end
always @(notifier_enable_h or notifier_slow)
begin
    disable LATCH_slow; slow_final <= 1'bx;
end
always @(*)
begin : LATCH_hld_ovr
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        hld_ovr_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        hld_ovr_final 	<= 1'b0;
    end
    else if (hld_h_n_buf===1)
    begin
        hld_ovr_final 	<= (^hld_ovr_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : hld_ovr_buf;
    end
end
always @(notifier_enable_h or notifier_hld_ovr)
begin
    disable LATCH_hld_ovr; hld_ovr_final <= 1'bx;
end
always @(*)
begin : LATCH_oe_n
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && (^hld_h_n_buf===1'bx || (hld_h_n_buf===0 && hld_ovr_final===1'bx)|| (hld_h_n_buf===1 && hld_ovr_final===1'bx))))
    begin
        oe_n_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        oe_n_final 	<= 1'b1;
    end
    else if (hld_h_n_buf===1 || hld_ovr_final===1)
    begin
        oe_n_final  	<= (^oe_n_buf  === 1'bx  || !pwr_good_hold_ovr_mode) ? 1'bx   : oe_n_buf;
    end
end
always @(notifier_enable_h or notifier_oe_n)
begin
    disable LATCH_oe_n; oe_n_final <= 1'bx;
end
always @(*)
begin : LATCH_out
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && (^hld_h_n_buf===1'bx ||(hld_h_n_buf===0 &&  hld_ovr_final===1'bx)||(hld_h_n_buf===1 &&  hld_ovr_final===1'bx))))
    begin
        out_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        out_final 	<= 1'b1;
    end
    else if (hld_h_n_buf===1 || hld_ovr_final===1)
    begin
        out_final  	<= (^out_buf  === 1'bx  || !pwr_good_hold_ovr_mode) ? 1'bx   : out_buf;
    end
end
always @(notifier_enable_h or notifier_out)
begin
    disable LATCH_out; out_final <= 1'bx;
end
always @(*)
begin
    if (x_on_analog_en_vdda ===1 )
    begin
        analog_en_vdda <= 1'bx;
    end
    else if ( zero_on_analog_en_vdda ===1 )
    begin
        analog_en_vdda <= 1'b0;
    end
    else if (x_on_analog_en_vdda !==1 && zero_on_analog_en_vdda !==1)
    begin
        analog_en_vdda <= ANALOG_EN;
    end
    if (x_on_analog_en_vddio_q  ===1 )
    begin
        analog_en_vddio_q  <= 1'bx;
    end
    else if ( zero_on_analog_en_vddio_q ===1 )
    begin
        analog_en_vddio_q  <= 1'b0;
    end
    else if ( x_on_analog_en_vddio_q !==1 && zero_on_analog_en_vddio_q !==1)
    begin
        analog_en_vddio_q  <= ANALOG_EN;
    end
    if (x_on_analog_en_vswitch  ===1 )
    begin
        analog_en_vswitch  <= 1'bx;
    end
    else if ( zero_on_analog_en_vswitch ===1 )
    begin
        analog_en_vswitch  <= 1'b0;
    end
    else if (x_on_analog_en_vswitch !==1 && zero_on_analog_en_vswitch !==1)
    begin
        analog_en_vswitch  <= ANALOG_EN;
    end
    if ( (analog_en_vswitch ===1'bx && analog_en_vdda ===1'bx) || (analog_en_vswitch ===1'bx && analog_en_vddio_q ===1'bx) || (analog_en_vddio_q ===1'bx && analog_en_vdda ===1'bx ) )
    begin
        analog_en_final  <= 1'bx;
    end
    else if (analog_en_vdda ===1'bx && (analog_en_vddio_q ===1 ||analog_en_vswitch===1 ))
    begin
        analog_en_final  <= 1'bx;
    end
    else if (analog_en_vddio_q ===1'bx && (analog_en_vdda ===1 ||analog_en_vswitch===1 ))
    begin
        analog_en_final  <= 1'bx;
    end
    else if (analog_en_vswitch===1'bx && (analog_en_vdda ===1 || analog_en_vddio_q ===1 ))
    begin
        analog_en_final  <= 1'bx;
    end
    else if ((analog_en_vdda ===0 && analog_en_vddio_q ===0 )|| (analog_en_vdda ===0 && analog_en_vswitch===0 ) ||  (analog_en_vddio_q ===0 && analog_en_vswitch===0 ))
    begin
        analog_en_final  <=0;
    end
    else if (analog_en_vdda ===1 && analog_en_vddio_q ===1 &&  analog_en_vswitch ===1)
    begin
        analog_en_final  <=1;
    end
end
wire [2:0] amux_select = {ANALOG_SEL, ANALOG_POL, out_buf};
wire invalid_controls_amux = 	(analog_en_final===1'bx && inp_dis_final===1)
     || !pwr_good_amux
     || (analog_en_final===1 && ^amux_select[2:0] === 1'bx && inp_dis_final===1);
wire enable_pad_amuxbus_a = invalid_controls_amux  ? 1'bx : (amux_select===3'b001 || amux_select===3'b010) && (analog_en_final===1);
wire enable_pad_amuxbus_b = invalid_controls_amux  ? 1'bx : (amux_select===3'b101 || amux_select===3'b110) && (analog_en_final===1);
wire enable_pad_vssio_q   = invalid_controls_amux  ? 1'bx : (amux_select===3'b100 || amux_select===3'b000) && (analog_en_final===1);
wire enable_pad_vddio_q   = invalid_controls_amux  ? 1'bx : (amux_select===3'b011 || amux_select===3'b111) && (analog_en_final===1);
tranif1 pad_amuxbus_a 	(PAD, AMUXBUS_A, enable_pad_amuxbus_a);
tranif1 pad_amuxbus_b 	(PAD, AMUXBUS_B, enable_pad_amuxbus_b);
bufif1 pad_vddio_q	(PAD, VDDIO_Q,   enable_pad_vddio_q);
bufif1 pad_vssio_q   	(PAD, VSSIO_Q,   enable_pad_vssio_q);
reg dis_err_msgs;
integer msg_count_pad,msg_count_pad1,msg_count_pad2,msg_count_pad3,msg_count_pad4,msg_count_pad5,msg_count_pad6,msg_count_pad7,msg_count_pad8,msg_count_pad9,msg_count_pad10,msg_count_pad11,msg_count_pad12;
initial
begin
    dis_err_msgs = 1'b1;
    msg_count_pad  = 0;
    msg_count_pad1 = 0;
    msg_count_pad2 = 0;
    msg_count_pad3 = 0;
    msg_count_pad4 = 0;
    msg_count_pad5 = 0;
    msg_count_pad6 = 0;
    msg_count_pad7 = 0;
    msg_count_pad8 = 0;
    msg_count_pad9 = 0;
    msg_count_pad10 = 0;
    msg_count_pad11 = 0;
    msg_count_pad12  = 0;


    #1;
    dis_err_msgs = 1'b0;

end
wire #100 error_enable_vddio = (ENABLE_VDDIO===0 && ENABLE_H===1);
event event_error_enable_vddio;
always @(error_enable_vddio)
begin
    if (!dis_err_msgs)
    begin
        if (error_enable_vddio===1)
        begin
            msg_count_pad = msg_count_pad + 1;
            ->event_error_enable_vddio;
            if (msg_count_pad <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 :  Enable_h (= %b) and ENABLE_VDDIO (= %b) are complement of each \other. This is an illegal combination as ENABLE_VDDIO and ENABLE_H are the same input signals IN different power \domains %m", ENABLE_H, ENABLE_VDDIO, $stime);
            end
            else
                if (msg_count_pad == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vdda = ( VDDA===1 && VDDIO_Q !==1 && ENABLE_VDDA_H===1 );
event event_error_vdda;
always @(error_vdda)
begin
    if (!dis_err_msgs)
    begin
        if (error_vdda===1)
        begin
            msg_count_pad1 = msg_count_pad1 + 1;
            ->event_error_vdda;
            if (msg_count_pad1 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ENABLE_VDDA_H (= %b) cannot be 1 when VDDA (= %b) and VDDIO_Q (= %b) %m",ENABLE_VDDA_H, VDDA,VDDIO_Q,$stime);
            end
            else
                if (msg_count_pad1 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vdda2 = ( VDDA===1 && VDDIO_Q ===1 && VSWITCH !==1 && ENABLE_H===1 && hld_h_n_buf ===1  &&  VCCD===1 && ANALOG_EN ===1 );
event event_error_vdda2;
always @(error_vdda2)
begin
    if (!dis_err_msgs)
    begin
        if (error_vdda2===1)
        begin
            msg_count_pad2 = msg_count_pad2 + 1;
            ->event_error_vdda2;
            if (msg_count_pad2 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ANALOG_EN (= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b), ENABLE_H (= %b),hld_h_n_buf (= %b) and VCCD (= %b)   %m",ANALOG_EN,VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,$stime);
            end
            else
                if (msg_count_pad2 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vdda3 =  ( VDDA===1 && VDDIO_Q ===1 && VSWITCH !==1 && ENABLE_H===1 && hld_h_n_buf ===1  && VCCD !==1 );
event event_error_vdda3;
always @(error_vdda3)
begin
    if (!dis_err_msgs)
    begin
        if (error_vdda3===1)
        begin
            msg_count_pad3 = msg_count_pad3 + 1;
            ->event_error_vdda3;
            if (msg_count_pad3 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : VCCD (= %b) cannot be any value other than 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b), ENABLE_H (= %b) and hld_h_n_buf (= %b) %m",VCCD,VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,$stime);
            end
            else
                if (msg_count_pad3 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch1 =  (VDDA !==1 && VDDIO_Q !==1 && VSWITCH ===1 && (ENABLE_VSWITCH_H===1)) ;
event event_error_vswitch1;
always @(error_vswitch1)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch1===1)
        begin
            msg_count_pad4 = msg_count_pad4 + 1;
            ->event_error_vswitch1;
            if (msg_count_pad4 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ENABLE_VSWITCH_H (= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) & VSWITCH(= %b) %m",ENABLE_VSWITCH_H,VDDA,VDDIO_Q,VSWITCH,$stime);
            end
            else
                if (msg_count_pad4 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch2 =   (VDDA !==1 && VDDIO_Q !==1 && VSWITCH ===1 && VCCD===1 && ANALOG_EN===1);
event event_error_vswitch2;
always @(error_vswitch2)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch2===1)
        begin
            msg_count_pad5 = msg_count_pad5 + 1;
            ->event_error_vswitch2;
            if (msg_count_pad5 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ANALOG_EN (= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b)  & VCCD(= %b) %m",ANALOG_EN,VDDA,VDDIO_Q,VSWITCH,VCCD,$stime);
            end
            else
                if (msg_count_pad5 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch3 =   (VDDA ===1 && VDDIO_Q !==1 && VSWITCH ===1 && ENABLE_VSWITCH_H===1);
event event_error_vswitch3;
always @(error_vswitch3)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch3===1)
        begin
            msg_count_pad6 = msg_count_pad6 + 1;
            ->event_error_vswitch3;
            if (msg_count_pad6 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ENABLE_VSWITCH_H(= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) & VSWITCH(= %b) %m",ENABLE_VSWITCH_H,VDDA,VDDIO_Q,VSWITCH,$stime);
            end
            else
                if (msg_count_pad6 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch4 =  (VDDA !==1 && VDDIO_Q ===1 && VSWITCH ===1 && ENABLE_VSWITCH_H===1);
event event_error_vswitch4;
always @(error_vswitch4)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch4===1)
        begin
            msg_count_pad7 = msg_count_pad7 + 1;
            ->event_error_vswitch4;
            if (msg_count_pad7 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ENABLE_VSWITCH_H(= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) & VSWITCH(= %b) %m",ENABLE_VSWITCH_H,VDDA,VDDIO_Q,VSWITCH,$stime);
            end
            else
                if (msg_count_pad7 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch5 =  (VDDA !==1 && VDDIO_Q ===1 && VSWITCH ===1 && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD ===1 && ANALOG_EN===1);
event event_error_vswitch5;
always @(error_vswitch5)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch5===1)
        begin
            msg_count_pad8 = msg_count_pad8 + 1;
            ->event_error_vswitch5;
            if (msg_count_pad8 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ANALOG_EN(= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b),ENABLE_H (= %b),hld_h_n_buf (= %b) and VCCD (= %b) %m",ANALOG_EN,VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,$stime);
            end
            else
                if (msg_count_pad8 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vddio_q1 =  (VDDA !==1 && VDDIO_Q ===1 && VSWITCH !==1 && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD!==1);
event event_error_vddio_q1;
always @(error_vddio_q1)
begin
    if (!dis_err_msgs)
    begin
        if (error_vddio_q1===1)
        begin
            msg_count_pad9 = msg_count_pad9 + 1;
            ->event_error_vddio_q1;
            if (msg_count_pad9 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : VCCD(= %b) cannot be any value other than 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b),ENABLE_H (= %b) and hld_h_n_buf (= %b)  %m",VCCD,VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,$stime);
            end
            else
                if (msg_count_pad9 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vddio_q2 =  (VDDA !==1 && VDDIO_Q ===1 && VSWITCH !==1 && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD ===1 && ANALOG_EN===1);
event event_error_vddio_q2;
always @(error_vddio_q2)
begin
    if (!dis_err_msgs)
    begin
        if (error_vddio_q2===1)
        begin
            msg_count_pad10 = msg_count_pad10 + 1;
            ->event_error_vddio_q2;
            if (msg_count_pad10 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ANALOG_EN(= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b),ENABLE_H (= %b) , hld_h_n_buf (= %b) && VCCD (= %b) %m",ANALOG_EN, VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,$stime);
            end
            else
                if (msg_count_pad10 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_supply_good = ( VDDA ===1 && VDDIO_Q ===1 && VSWITCH ===1  && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD ===1 &&  ANALOG_EN===1 && ENABLE_VSWITCH_H !==1 && ENABLE_VSWITCH_H !==0 );
event event_error_supply_good;
always @(error_supply_good)
begin
    if (!dis_err_msgs)
    begin
        if (error_supply_good===1)
        begin
            msg_count_pad11 = msg_count_pad11 + 1;
            ->event_error_supply_good;
            if (msg_count_pad11 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ENABLE_VSWITCH_H(= %b) should be either 1 or 0 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b), ENABLE_H (= %b), hld_h_n_buf (= %b) ,VCCD (= %b) and ANALOG_EN(= %b)  %m",ENABLE_VSWITCH_H, VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,ANALOG_EN,$stime);
            end
            else
                if (msg_count_pad11 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vdda_vddioq_vswitch2 = ( VDDA ===1 && VDDIO_Q ===1 && VSWITCH ===1 && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD ===1 &&  ANALOG_EN===1 && ENABLE_VDDA_H !==1 && ENABLE_VDDA_H !==0 );
event event_error_vdda_vddioq_vswitch2;
always @(error_vdda_vddioq_vswitch2)
begin
    if (!dis_err_msgs)
    begin
        if (error_vdda_vddioq_vswitch2===1)
        begin
            msg_count_pad12 = msg_count_pad12 + 1;
            ->event_error_vdda_vddioq_vswitch2;
            if (msg_count_pad12 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpio_ovtv2 : ENABLE_VDDA_H(= %b) should be either 1 or 0 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b), ENABLE_H (= %b), hld_h_n_buf (= %b) ,VCCD (= %b) and ANALOG_EN(= %b)  %m",ENABLE_VDDA_H, VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,ANALOG_EN,$stime);
            end
            else
                if (msg_count_pad12 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpio_ovtv2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
endmodule


















































































































































































































































































































































































































































































































































































































































































































































































































































































































































 // FUNCTIONAL















































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_GPIO_OVTV2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_gpiov2: General Purpose I/0.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_gpiov2 (IN_H, PAD_A_NOESD_H,PAD_A_ESD_0_H,PAD_A_ESD_1_H,
                                 PAD, DM, HLD_H_N, IN, INP_DIS, IB_MODE_SEL, ENABLE_H, ENABLE_VDDA_H, ENABLE_INP_H, OE_N,
                                 TIE_HI_ESD, TIE_LO_ESD, SLOW, VTRIP_SEL, HLD_OVR, ANALOG_EN, ANALOG_SEL, ENABLE_VDDIO, ENABLE_VSWITCH_H,
                                 ANALOG_POL, OUT, AMUXBUS_A, AMUXBUS_B
                                 ,VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VSSIO,
                                 VSSD, VSSIO_Q
                                );
input OUT;
input OE_N;
input HLD_H_N;
input ENABLE_H;
input ENABLE_INP_H;
input ENABLE_VDDA_H;
input ENABLE_VSWITCH_H;
input ENABLE_VDDIO;
input INP_DIS;
input IB_MODE_SEL;
input VTRIP_SEL;
input SLOW;
input HLD_OVR;
input ANALOG_EN;
input ANALOG_SEL;
input ANALOG_POL;
input [2:0] DM;
inout VDDIO;
inout VDDIO_Q;
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;
inout PAD;
inout PAD_A_NOESD_H,PAD_A_ESD_0_H,PAD_A_ESD_1_H;
inout AMUXBUS_A;
inout AMUXBUS_B;
output IN;
output IN_H;
output TIE_HI_ESD, TIE_LO_ESD;
reg [2:0] dm_final;
reg slow_final, vtrip_sel_final, inp_dis_final, out_final, oe_n_final, hld_ovr_final, analog_en_final, ib_mode_sel_final, analog_en_vdda, analog_en_vswitch,analog_en_vddio_q;
wire [2:0] dm_buf;
wire slow_buf, vtrip_sel_buf, inp_dis_buf, out_buf, oe_n_buf, hld_ovr_buf,ib_mode_sel_buf;
wire [2:0] dm_del;
wire slow_del, vtrip_sel_del, inp_dis_del, out_del, oe_n_del, hld_ovr_del,ib_mode_sel_del;
wire hld_h_n_del;
wire hld_h_n_buf;
reg notifier_dm, notifier_slow, notifier_oe_n, notifier_out, notifier_vtrip_sel, notifier_hld_ovr, notifier_inp_dis, notifier_ib_mode_sel;
reg notifier_enable_h, notifier;
assign hld_h_n_buf 	= HLD_H_N;
assign hld_ovr_buf 	= HLD_OVR;
assign dm_buf 		= DM;
assign inp_dis_buf 	= INP_DIS;
assign vtrip_sel_buf 	= VTRIP_SEL;
assign slow_buf 	= SLOW;
assign oe_n_buf 	= OE_N;
assign out_buf 		= OUT;
assign ib_mode_sel_buf 	= IB_MODE_SEL;
wire  pwr_good_amux	       = ((hld_h_n_buf===0 || ENABLE_H===0) ? 1:(VCCD===1))  && (VSSD===0) && (VSSA===0) && (VSSIO_Q===0);
wire  pwr_good_hold_ovr_mode   = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0)    && (VCCHIB===1);
wire  pwr_good_active_mode     = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0)    && (VCCD===1);
wire  pwr_good_hold_mode       = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0);
wire  pwr_good_active_mode_vdda = (VDDA===1)  && (VSSD===0)   && (VCCD===1);
wire  pwr_good_hold_mode_vdda   = (VDDA===1)    && (VSSD===0);
wire  pwr_good_inpbuff_hv       = (VDDIO_Q===1) && (VSSD===0)   && (inp_dis_final===0 && dm_final!==3'b000 && ib_mode_sel_final===1 ? VCCHIB===1 : 1);
wire  pwr_good_inpbuff_lv       = (VDDIO_Q===1) && (VSSD===0)   && (VCCHIB===1);
wire  pwr_good_output_driver    = (VDDIO===1)   && (VDDIO_Q===1)&& (VSSIO===0)   && (VSSD===0)  && (VSSA===0) ;
wire  pwr_good_analog_en_vdda   = (VDDA===1)  && (VSSD===0) && (VSSA===0) ;
wire  pwr_good_analog_en_vddio_q = (VDDIO_Q ===1)  && (VSSD===0) && (VSSA===0) ;
wire  pwr_good_analog_en_vswitch = (VSWITCH ===1)  && (VSSD===0) && (VSSA===0) ;
wire  pwr_good_amux_vccd   = ((hld_h_n_buf===0 || ENABLE_H===0) ? 1:(VCCD===1));
parameter MAX_WARNING_COUNT = 100;
wire pad_tristate = oe_n_final === 1 || dm_final === 3'b000 || dm_final === 3'b001;
wire x_on_pad  =  !pwr_good_output_driver
     || (dm_final !== 3'b000 && dm_final !== 3'b001 && oe_n_final===1'bx)
     || (^dm_final[2:0] === 1'bx && oe_n_final===1'b0)
     || (slow_final===1'bx && dm_final !== 3'b000 && dm_final !== 3'b001 && oe_n_final===1'b0);




parameter SLOW_1_DELAY= 0;
parameter SLOW_0_DELAY= 0;

integer slow_1_delay,slow_0_delay,slow_delay;
initial slow_1_delay = SLOW_1_DELAY;
initial slow_0_delay = SLOW_0_DELAY;
always @(*)
begin
    if (SLOW===1)
        slow_delay = slow_1_delay;
    else
        slow_delay = slow_0_delay;
end
bufif1 (pull1, strong0) #slow_delay dm2 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b010));
bufif1 (strong1, pull0) #slow_delay dm3 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b011));
bufif1 (highz1, strong0) #slow_delay dm4 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b100));
bufif1 (strong1, highz0) #slow_delay dm5 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b101));
bufif1 (strong1, strong0) #slow_delay dm6 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b110));
bufif1 (pull1, pull0)  #slow_delay dm7 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b111));
tran pad_esd_1 (PAD,PAD_A_NOESD_H);
tran pad_esd_2 (PAD,PAD_A_ESD_0_H);
tran pad_esd_3 (PAD,PAD_A_ESD_1_H);
wire x_on_in_hv  =  (ENABLE_H===0  && ^ENABLE_INP_H===1'bx)
     || (inp_dis_final===1'bx  && ^dm_final[2:0]!==1'bx && dm_final !== 3'b000)
     || (^ENABLE_H===1'bx)
     || (inp_dis_final===0 	       	&& ^dm_final[2:0] === 1'bx)
     || (ib_mode_sel_final===1'bx  	&& inp_dis_final===0        && dm_final !== 3'b000)
     || (^ENABLE_VDDIO===1'bx    	&& inp_dis_final===0        && dm_final !== 3'b000	&& ib_mode_sel_final===1'b1)
     || (vtrip_sel_final===1'bx    	&& inp_dis_final===0        && dm_final !== 3'b000	&& ib_mode_sel_final===1'b0);
wire x_on_in_lv  =  (ENABLE_H===0  && ^ENABLE_INP_H===1'bx)
     || (inp_dis_final===1'bx  && ^dm_final[2:0]!==1'bx && dm_final !== 3'b000)
     || (ENABLE_H===0  && ^ENABLE_VDDIO===1'bx)
     || (^ENABLE_H===1'bx)
     || (inp_dis_final===0 	       	&& ^dm_final[2:0] === 1'bx)
     || (ib_mode_sel_final===1'bx  	&& inp_dis_final===0        && dm_final !== 3'b000)
     || (^ENABLE_VDDIO===1'bx    	&& inp_dis_final===0        && dm_final !== 3'b000)
     || (vtrip_sel_final===1'bx    	&& inp_dis_final===0        && dm_final !== 3'b000	&& ib_mode_sel_final===1'b0);
wire disable_inp_buff = ENABLE_H===1 ? (dm_final===3'b000 || inp_dis_final===1) : ENABLE_INP_H===0;
assign IN_H = (x_on_in_hv===1 || pwr_good_inpbuff_hv===0) ? 1'bx : (disable_inp_buff===1 ? 0 : (^PAD===1'bx ? 1'bx : PAD));
wire disable_inp_buff_lv = ENABLE_H===1 ? (dm_final===3'b000 || inp_dis_final===1) : ENABLE_VDDIO===0;
assign IN =   (x_on_in_lv===1 || pwr_good_inpbuff_lv===0 ) ? 1'bx : (disable_inp_buff_lv===1 ? 0 : (^PAD===1'bx ? 1'bx : PAD));
assign TIE_HI_ESD = VDDIO===1'b1 ? 1'b1 : 1'bx;
assign TIE_LO_ESD = VSSIO===1'b0 ? 1'b0 : 1'bx;
wire functional_mode_amux = (pwr_good_analog_en_vdda ===1 && pwr_good_analog_en_vddio_q ===1 && pwr_good_analog_en_vswitch ===1 );
wire x_on_analog_en_vdda = (pwr_good_analog_en_vdda !==1
                            || (functional_mode_amux ==1 && (ENABLE_H !==0 && ^hld_h_n_buf === 1'bx) || (hld_h_n_buf!== 0 && ^ENABLE_H=== 1'bx) || pwr_good_amux_vccd !==1 )
                            || (functional_mode_amux ==1 && (hld_h_n_buf ===1 && ENABLE_H===1 && ^ANALOG_EN === 1'bx && ENABLE_VDDA_H ===1 && ENABLE_VSWITCH_H===1 ) || (hld_h_n_buf ===1 && ENABLE_H===1 && ANALOG_EN ===0 && ^ENABLE_VDDA_H ===1'bx) ));
wire zero_on_analog_en_vdda = ( (pwr_good_analog_en_vdda ===1 && ENABLE_VDDA_H ===0)
                                || (pwr_good_analog_en_vdda ===1 && pwr_good_analog_en_vddio_q ===1 && hld_h_n_buf===0)
                                || (pwr_good_analog_en_vdda ===1 && pwr_good_analog_en_vddio_q ===1 && ENABLE_H===0)
                                ||  (pwr_good_analog_en_vdda ===1 && pwr_good_analog_en_vddio_q ===1 && pwr_good_amux_vccd && ANALOG_EN===0) );
wire x_on_analog_en_vddio_q =  ( pwr_good_analog_en_vddio_q !==1
                                 || (functional_mode_amux ==1 && (ENABLE_H !==0 && ^hld_h_n_buf === 1'bx) || (hld_h_n_buf!== 0 && ^ENABLE_H=== 1'bx) || pwr_good_amux_vccd !==1 )
                                 || (functional_mode_amux ==1 && (hld_h_n_buf ===1 && ENABLE_H===1 && ^ANALOG_EN === 1'bx && ENABLE_VDDA_H ===1 && ENABLE_VSWITCH_H===1 ) ));
wire zero_on_analog_en_vddio_q =  ( (pwr_good_analog_en_vddio_q ===1 && hld_h_n_buf===0)
                                    || (pwr_good_analog_en_vddio_q ===1 && ENABLE_H===0)
                                    ||  (pwr_good_analog_en_vddio_q ===1 && pwr_good_amux_vccd && ANALOG_EN===0) );
wire x_on_analog_en_vswitch = (pwr_good_analog_en_vswitch !==1
                               || (functional_mode_amux ==1 && (ENABLE_H !==0 && ^hld_h_n_buf === 1'bx) || (hld_h_n_buf!== 0 && ^ENABLE_H=== 1'bx) || pwr_good_amux_vccd !==1 )
                               || (functional_mode_amux ==1 && (hld_h_n_buf ===1 && ENABLE_H===1 && ^ANALOG_EN === 1'bx && ENABLE_VDDA_H ===1 && ENABLE_VSWITCH_H===1 ) || (hld_h_n_buf ===1 && ENABLE_H===1 && ANALOG_EN ===0 && ^ENABLE_VSWITCH_H ===1'bx) ));
wire  zero_on_analog_en_vswitch =   ( (pwr_good_analog_en_vswitch ===1 && ENABLE_VSWITCH_H ===0)
                                      || (pwr_good_analog_en_vswitch ===1 && pwr_good_analog_en_vddio_q ===1 && hld_h_n_buf===0)
                                      || (pwr_good_analog_en_vswitch ===1 && pwr_good_analog_en_vddio_q ===1 && ENABLE_H===0)
                                      ||  (pwr_good_analog_en_vswitch ===1 && pwr_good_analog_en_vddio_q ===1 && pwr_good_amux_vccd && ANALOG_EN===0) );
always @(*)
begin : LATCH_dm
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        dm_final 	<= 3'bxxx;
    end
    else if (ENABLE_H===0)
    begin
        dm_final 	<= 3'b000;
    end
    else if (hld_h_n_buf===1)
    begin
        dm_final 	<= (^dm_buf[2:0]	=== 1'bx	|| !pwr_good_active_mode) ? 3'bxxx : dm_buf;
    end
end
always @(notifier_enable_h or notifier_dm)
begin
    disable LATCH_dm; dm_final <= 3'bxxx;
end
always @(*)
begin : LATCH_inp_dis
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        inp_dis_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        inp_dis_final 	<= 1'b1;
    end
    else if (hld_h_n_buf===1)
    begin
        inp_dis_final 	<= (^inp_dis_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : inp_dis_buf;
    end
end
always @(notifier_enable_h or notifier_inp_dis)
begin
    disable LATCH_inp_dis; inp_dis_final <= 1'bx;
end
always @(*)
begin : LATCH_vtrip_sel
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        vtrip_sel_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        vtrip_sel_final 	<= 1'b0;
    end
    else if (hld_h_n_buf===1)
    begin
        vtrip_sel_final 	<= (^vtrip_sel_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : vtrip_sel_buf;
    end
end
always @(notifier_enable_h or notifier_vtrip_sel)
begin
    disable LATCH_vtrip_sel; vtrip_sel_final <= 1'bx;
end
always @(*)
begin : LATCH_ib_mode_sel
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        ib_mode_sel_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        ib_mode_sel_final 	<= 1'b0;
    end
    else if (hld_h_n_buf===1)
    begin
        ib_mode_sel_final 	<= (^ib_mode_sel_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : ib_mode_sel_buf;
    end
end
always @(notifier_enable_h or notifier_ib_mode_sel)
begin
    disable LATCH_ib_mode_sel; ib_mode_sel_final <= 1'bx;
end
always @(*)
begin : LATCH_slow
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        slow_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        slow_final 	<= 1'b0;
    end
    else if (hld_h_n_buf===1)
    begin
        slow_final 	<= (^slow_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : slow_buf;
    end
end
always @(notifier_enable_h or notifier_slow)
begin
    disable LATCH_slow; slow_final <= 1'bx;
end
always @(*)
begin : LATCH_hld_ovr
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^hld_h_n_buf===1'bx))
    begin
        hld_ovr_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        hld_ovr_final 	<= 1'b0;
    end
    else if (hld_h_n_buf===1)
    begin
        hld_ovr_final 	<= (^hld_ovr_buf === 1'bx	|| !pwr_good_active_mode) ? 1'bx : hld_ovr_buf;
    end
end
always @(notifier_enable_h or notifier_hld_ovr)
begin
    disable LATCH_hld_ovr; hld_ovr_final <= 1'bx;
end
always @(*)
begin : LATCH_oe_n
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && (^hld_h_n_buf===1'bx || (hld_h_n_buf===0 && hld_ovr_final===1'bx) || (hld_h_n_buf===1 && hld_ovr_final===1'bx))))
    begin
        oe_n_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        oe_n_final 	<= 1'b1;
    end
    else if (hld_h_n_buf===1 || hld_ovr_final===1)
    begin
        oe_n_final  	<= (^oe_n_buf  === 1'bx  || !pwr_good_hold_ovr_mode) ? 1'bx   : oe_n_buf;
    end
end
always @(notifier_enable_h or notifier_oe_n)
begin
    disable LATCH_oe_n; oe_n_final <= 1'bx;
end
always @(*)
begin : LATCH_out
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && (^hld_h_n_buf===1'bx ||(hld_h_n_buf===0 &&  hld_ovr_final===1'bx || (hld_h_n_buf===1 && hld_ovr_final===1'bx)))))
    begin
        out_final 	<= 1'bx;
    end
    else if (ENABLE_H===0)
    begin
        out_final 	<= 1'b1;
    end
    else if (hld_h_n_buf===1 || hld_ovr_final===1)
    begin
        out_final  	<= (^out_buf  === 1'bx  || !pwr_good_hold_ovr_mode) ? 1'bx   : out_buf;
    end
end
always @(notifier_enable_h or notifier_out)
begin
    disable LATCH_out; out_final <= 1'bx;
end
always @(*)
begin
    if (x_on_analog_en_vdda ===1 )
    begin
        analog_en_vdda <= 1'bx;
    end
    else if ( zero_on_analog_en_vdda ===1 )
    begin
        analog_en_vdda <= 1'b0;
    end
    else if (x_on_analog_en_vdda !==1 && zero_on_analog_en_vdda !==1)
    begin
        analog_en_vdda <= ANALOG_EN;
    end
    if (x_on_analog_en_vddio_q  ===1 )
    begin
        analog_en_vddio_q  <= 1'bx;
    end
    else if ( zero_on_analog_en_vddio_q ===1 )
    begin
        analog_en_vddio_q  <= 1'b0;
    end
    else if ( x_on_analog_en_vddio_q !==1 && zero_on_analog_en_vddio_q !==1)
    begin
        analog_en_vddio_q  <= ANALOG_EN;
    end
    if (x_on_analog_en_vswitch  ===1 )
    begin
        analog_en_vswitch  <= 1'bx;
    end
    else if ( zero_on_analog_en_vswitch ===1 )
    begin
        analog_en_vswitch  <= 1'b0;
    end
    else if (x_on_analog_en_vswitch !==1 && zero_on_analog_en_vswitch !==1)
    begin
        analog_en_vswitch  <= ANALOG_EN;
    end
    if ( (analog_en_vswitch ===1'bx && analog_en_vdda ===1'bx) || (analog_en_vswitch ===1'bx && analog_en_vddio_q ===1'bx) || (analog_en_vddio_q ===1'bx && analog_en_vdda ===1'bx ) )
    begin
        analog_en_final  <= 1'bx;
    end
    else if (analog_en_vdda ===1'bx && (analog_en_vddio_q ===1 ||analog_en_vswitch===1 ))
    begin
        analog_en_final  <= 1'bx;
    end
    else if (analog_en_vddio_q ===1'bx && (analog_en_vdda ===1 ||analog_en_vswitch===1 ))
    begin
        analog_en_final  <= 1'bx;
    end
    else if (analog_en_vswitch===1'bx && (analog_en_vdda ===1 || analog_en_vddio_q ===1 ))
    begin
        analog_en_final  <= 1'bx;
    end
    else if ((analog_en_vdda ===0 && analog_en_vddio_q ===0 )|| (analog_en_vdda ===0 && analog_en_vswitch===0 ) ||  (analog_en_vddio_q ===0 && analog_en_vswitch===0 ))
    begin
        analog_en_final  <=0;
    end
    else if (analog_en_vdda ===1 && analog_en_vddio_q ===1 &&  analog_en_vswitch ===1)
    begin
        analog_en_final  <=1;
    end
end
wire [2:0] amux_select = {ANALOG_SEL, ANALOG_POL, out_buf};
wire invalid_controls_amux = 	(analog_en_final===1'bx && inp_dis_final===1)
     || !pwr_good_amux
     || (analog_en_final===1 && ^amux_select[2:0] === 1'bx && inp_dis_final===1);
wire enable_pad_amuxbus_a = invalid_controls_amux  ? 1'bx : (amux_select===3'b001 || amux_select===3'b010) && (analog_en_final===1);
wire enable_pad_amuxbus_b = invalid_controls_amux  ? 1'bx : (amux_select===3'b101 || amux_select===3'b110) && (analog_en_final===1);
wire enable_pad_vssio_q   = invalid_controls_amux  ? 1'bx : (amux_select===3'b100 || amux_select===3'b000) && (analog_en_final===1);
wire enable_pad_vddio_q   = invalid_controls_amux  ? 1'bx : (amux_select===3'b011 || amux_select===3'b111) && (analog_en_final===1);
tranif1 pad_amuxbus_a 	(PAD, AMUXBUS_A, enable_pad_amuxbus_a);
tranif1 pad_amuxbus_b 	(PAD, AMUXBUS_B, enable_pad_amuxbus_b);
bufif1 pad_vddio_q	(PAD, VDDIO_Q,   enable_pad_vddio_q);
bufif1 pad_vssio_q   	(PAD, VSSIO_Q,   enable_pad_vssio_q);
reg dis_err_msgs;
integer msg_count_pad,msg_count_pad1,msg_count_pad2,msg_count_pad3,msg_count_pad4,msg_count_pad5,msg_count_pad6,msg_count_pad7,msg_count_pad8,msg_count_pad9,msg_count_pad10,msg_count_pad11,msg_count_pad12;
initial
begin
    dis_err_msgs = 1'b1;
    msg_count_pad  = 0;
    msg_count_pad1 = 0;
    msg_count_pad2 = 0;
    msg_count_pad3 = 0;
    msg_count_pad4 = 0;
    msg_count_pad5 = 0;
    msg_count_pad6 = 0;
    msg_count_pad7 = 0;
    msg_count_pad8 = 0;
    msg_count_pad9 = 0;
    msg_count_pad10 = 0;
    msg_count_pad11 = 0;
    msg_count_pad12  = 0;


    #1;
    dis_err_msgs = 1'b0;

end
wire #100 error_enable_vddio = (ENABLE_VDDIO===0 && ENABLE_H===1);
event event_error_enable_vddio;
always @(error_enable_vddio)
begin
    if (!dis_err_msgs)
    begin
        if (error_enable_vddio===1)
        begin
            msg_count_pad = msg_count_pad + 1;
            ->event_error_enable_vddio;
            if (msg_count_pad <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 :  Enable_h (= %b) and ENABLE_VDDIO (= %b) are complement of each \other. This is an illegal combination as ENABLE_VDDIO and ENABLE_H are the same input signals IN different power \domains %m", ENABLE_H, ENABLE_VDDIO, $stime);
            end
            else
                if (msg_count_pad == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vdda = ( VDDA===1 && VDDIO_Q !==1 && ENABLE_VDDA_H===1 );
event event_error_vdda;
always @(error_vdda)
begin
    if (!dis_err_msgs)
    begin
        if (error_vdda===1)
        begin
            msg_count_pad1 = msg_count_pad1 + 1;
            ->event_error_vdda;
            if (msg_count_pad1 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ENABLE_VDDA_H (= %b) cannot be 1 when VDDA (= %b) and VDDIO_Q (= %b) %m",ENABLE_VDDA_H, VDDA,VDDIO_Q,$stime);
            end
            else
                if (msg_count_pad1 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vdda2 = ( VDDA===1 && VDDIO_Q ===1 && VSWITCH !==1 && ENABLE_H===1 && hld_h_n_buf ===1  &&  VCCD===1 && ANALOG_EN ===1 );
event event_error_vdda2;
always @(error_vdda2)
begin
    if (!dis_err_msgs)
    begin
        if (error_vdda2===1)
        begin
            msg_count_pad2 = msg_count_pad2 + 1;
            ->event_error_vdda2;
            if (msg_count_pad2 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ANALOG_EN (= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b), ENABLE_H (= %b),hld_h_n_buf (= %b) and VCCD (= %b)   %m",ANALOG_EN,VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,$stime);
            end
            else
                if (msg_count_pad2 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vdda3 =  ( VDDA===1 && VDDIO_Q ===1 && VSWITCH !==1 && ENABLE_H===1 && hld_h_n_buf ===1  && VCCD !==1 );
event event_error_vdda3;
always @(error_vdda3)
begin
    if (!dis_err_msgs)
    begin
        if (error_vdda3===1)
        begin
            msg_count_pad3 = msg_count_pad3 + 1;
            ->event_error_vdda3;
            if (msg_count_pad3 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : VCCD (= %b) cannot be any value other than 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b), ENABLE_H (= %b) and hld_h_n_buf (= %b) %m",VCCD,VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,$stime);
            end
            else
                if (msg_count_pad3 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch1 =  (VDDA !==1 && VDDIO_Q !==1 && VSWITCH ===1 && (ENABLE_VSWITCH_H===1)) ;
event event_error_vswitch1;
always @(error_vswitch1)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch1===1)
        begin
            msg_count_pad4 = msg_count_pad4 + 1;
            ->event_error_vswitch1;
            if (msg_count_pad4 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ENABLE_VSWITCH_H (= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) & VSWITCH(= %b) %m",ENABLE_VSWITCH_H,VDDA,VDDIO_Q,VSWITCH,$stime);
            end
            else
                if (msg_count_pad4 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch2 =   (VDDA !==1 && VDDIO_Q !==1 && VSWITCH ===1 && VCCD===1 && ANALOG_EN===1);
event event_error_vswitch2;
always @(error_vswitch2)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch2===1)
        begin
            msg_count_pad5 = msg_count_pad5 + 1;
            ->event_error_vswitch2;
            if (msg_count_pad5 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ANALOG_EN (= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b)  & VCCD(= %b) %m",ANALOG_EN,VDDA,VDDIO_Q,VSWITCH,VCCD,$stime);
            end
            else
                if (msg_count_pad5 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch3 =   (VDDA ===1 && VDDIO_Q !==1 && VSWITCH ===1 && ENABLE_VSWITCH_H===1);
event event_error_vswitch3;
always @(error_vswitch3)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch3===1)
        begin
            msg_count_pad6 = msg_count_pad6 + 1;
            ->event_error_vswitch3;
            if (msg_count_pad6 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ENABLE_VSWITCH_H(= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) & VSWITCH(= %b) %m",ENABLE_VSWITCH_H,VDDA,VDDIO_Q,VSWITCH,$stime);
            end
            else
                if (msg_count_pad6 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch4 =  (VDDA !==1 && VDDIO_Q ===1 && VSWITCH ===1 && ENABLE_VSWITCH_H===1);
event event_error_vswitch4;
always @(error_vswitch4)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch4===1)
        begin
            msg_count_pad7 = msg_count_pad7 + 1;
            ->event_error_vswitch4;
            if (msg_count_pad7 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ENABLE_VSWITCH_H(= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) & VSWITCH(= %b) %m",ENABLE_VSWITCH_H,VDDA,VDDIO_Q,VSWITCH,$stime);
            end
            else
                if (msg_count_pad7 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vswitch5 =  (VDDA !==1 && VDDIO_Q ===1 && VSWITCH ===1 && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD ===1 && ANALOG_EN===1);
event event_error_vswitch5;
always @(error_vswitch5)
begin
    if (!dis_err_msgs)
    begin
        if (error_vswitch5===1)
        begin
            msg_count_pad8 = msg_count_pad8 + 1;
            ->event_error_vswitch5;
            if (msg_count_pad8 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ANALOG_EN(= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b),ENABLE_H (= %b),hld_h_n_buf (= %b) and VCCD (= %b) %m",ANALOG_EN,VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,$stime);
            end
            else
                if (msg_count_pad8 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vddio_q1 =  (VDDA !==1 && VDDIO_Q ===1 && VSWITCH !==1 && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD!==1);
event event_error_vddio_q1;
always @(error_vddio_q1)
begin
    if (!dis_err_msgs)
    begin
        if (error_vddio_q1===1)
        begin
            msg_count_pad9 = msg_count_pad9 + 1;
            ->event_error_vddio_q1;
            if (msg_count_pad9 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : VCCD(= %b) cannot be any value other than 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b),ENABLE_H (= %b) and hld_h_n_buf (= %b)  %m",VCCD,VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,$stime);
            end
            else
                if (msg_count_pad9 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vddio_q2 =  (VDDA !==1 && VDDIO_Q ===1 && VSWITCH !==1 && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD ===1 && ANALOG_EN===1);
event event_error_vddio_q2;
always @(error_vddio_q2)
begin
    if (!dis_err_msgs)
    begin
        if (error_vddio_q2===1)
        begin
            msg_count_pad10 = msg_count_pad10 + 1;
            ->event_error_vddio_q2;
            if (msg_count_pad10 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ANALOG_EN(= %b) cannot be 1 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b),ENABLE_H (= %b) , hld_h_n_buf (= %b) && VCCD (= %b) %m",ANALOG_EN, VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,$stime);
            end
            else
                if (msg_count_pad10 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_supply_good = ( VDDA ===1 && VDDIO_Q ===1 && VSWITCH ===1  && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD ===1 &&  ANALOG_EN===1 && ENABLE_VSWITCH_H !==1 && ENABLE_VSWITCH_H !==0 );
event event_error_supply_good;
always @(error_supply_good)
begin
    if (!dis_err_msgs)
    begin
        if (error_supply_good===1)
        begin
            msg_count_pad11 = msg_count_pad11 + 1;
            ->event_error_supply_good;
            if (msg_count_pad11 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ENABLE_VSWITCH_H(= %b) should be either 1 or 0 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b), ENABLE_H (= %b), hld_h_n_buf (= %b) ,VCCD (= %b) and ANALOG_EN(= %b)  %m",ENABLE_VSWITCH_H, VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,ANALOG_EN,$stime);
            end
            else
                if (msg_count_pad11 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
wire #100 error_vdda_vddioq_vswitch2 = ( VDDA ===1 && VDDIO_Q ===1 && VSWITCH ===1 && ENABLE_H ===1 && hld_h_n_buf ===1 && VCCD ===1 &&  ANALOG_EN===1 && ENABLE_VDDA_H !==1 && ENABLE_VDDA_H !==0 );
event event_error_vdda_vddioq_vswitch2;
always @(error_vdda_vddioq_vswitch2)
begin
    if (!dis_err_msgs)
    begin
        if (error_vdda_vddioq_vswitch2===1)
        begin
            msg_count_pad12 = msg_count_pad12 + 1;
            ->event_error_vdda_vddioq_vswitch2;
            if (msg_count_pad12 <= MAX_WARNING_COUNT)
            begin
                $display(" ===ERROR=== sky130_fd_io__top_gpiov2 : ENABLE_VDDA_H(= %b) should be either 1 or 0 when VDDA (= %b) , VDDIO_Q (= %b) , VSWITCH(= %b), ENABLE_H (= %b), hld_h_n_buf (= %b) ,VCCD (= %b) and ANALOG_EN(= %b)  %m",ENABLE_VDDA_H, VDDA,VDDIO_Q,VSWITCH,ENABLE_H,hld_h_n_buf,VCCD,ANALOG_EN,$stime);
            end
            else
                if (msg_count_pad12 == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_gpiov2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
endmodule






























































































































































































































































































































































































































































































































































































































































































































































































































 // FUNCTIONAL



































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_GPIOV2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_ground_hvc_wpad: Ground pad.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_ground_hvc_wpad ( G_PAD, AMUXBUS_A, AMUXBUS_B
        , G_CORE, DRN_HVC, OGC_HVC, SRC_BDY_HVC,VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VSSIO, VSSD, VSSIO_Q
                                         );
inout G_PAD;
inout AMUXBUS_A;
inout AMUXBUS_B;
inout OGC_HVC;
inout DRN_HVC;
inout SRC_BDY_HVC;
inout G_CORE;
inout VDDIO;
inout VDDIO_Q;
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;
assign G_CORE = G_PAD;
endmodule









































 // FUNCTIONAL

























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_GROUND_HVC_WPAD_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_ground_lvc_wpad: Base ground I/O pad with low voltage clamp.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_ground_lvc_wpad ( G_PAD, AMUXBUS_A, AMUXBUS_B
        , G_CORE, BDY2_B2B, DRN_LVC1, DRN_LVC2, OGC_LVC, SRC_BDY_LVC1, SRC_BDY_LVC2, VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VSSIO, VSSD, VSSIO_Q
                                         );
inout G_PAD;
inout AMUXBUS_A;
inout AMUXBUS_B;
inout SRC_BDY_LVC1;
inout SRC_BDY_LVC2;
inout OGC_LVC;
inout DRN_LVC1;
inout BDY2_B2B;
inout DRN_LVC2;
inout G_CORE;
inout VDDIO;
inout VDDIO_Q;
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;
assign G_CORE = G_PAD;
endmodule












































 // FUNCTIONAL































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_GROUND_LVC_WPAD_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_power_hvc_wpad: A power pad with an ESD high-voltage clamp.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_power_hvc_wpad ( P_PAD, AMUXBUS_A, AMUXBUS_B
        , P_CORE, DRN_HVC, OGC_HVC, SRC_BDY_HVC,VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VSSIO, VSSD, VSSIO_Q
                                        );
inout P_PAD;
inout AMUXBUS_A;
inout AMUXBUS_B;
inout OGC_HVC;
inout DRN_HVC;
inout SRC_BDY_HVC;
inout P_CORE;
inout VDDIO;
inout VDDIO_Q;
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;
assign P_CORE = P_PAD;
endmodule









































 // FUNCTIONAL

























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_POWER_HVC_WPAD_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_power_hvc_wpadv2: A power pad with an ESD high-voltage clamp.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_power_hvc_wpadv2 ( P_PAD, AMUXBUS_A, AMUXBUS_B
        , P_CORE, DRN_HVC, OGC_HVC, SRC_BDY_HVC,VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VSSIO, VSSD, VSSIO_Q
                                          );
inout P_PAD;
inout AMUXBUS_A;
inout AMUXBUS_B;
inout OGC_HVC;
inout DRN_HVC;
inout SRC_BDY_HVC;
inout P_CORE;
inout VDDIO;
inout VDDIO_Q;
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;
tran p1 (P_CORE, P_PAD);
endmodule









































 // FUNCTIONAL

























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_POWER_HVC_WPADV2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_power_lvc_wpad: A power pad with an ESD low-voltage clamp.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_power_lvc_wpad ( P_PAD, AMUXBUS_A, AMUXBUS_B
        , P_CORE, BDY2_B2B, DRN_LVC1, DRN_LVC2, OGC_LVC, SRC_BDY_LVC1, SRC_BDY_LVC2, VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VSSIO, VSSD, VSSIO_Q
                                        );
inout P_PAD;
inout AMUXBUS_A;
inout AMUXBUS_B;
inout SRC_BDY_LVC1;
inout SRC_BDY_LVC2;
inout OGC_LVC;
inout DRN_LVC1;
inout BDY2_B2B;
inout DRN_LVC2;
inout P_CORE;
inout VDDIO;
inout VDDIO_Q;
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;
assign P_CORE = P_PAD;
endmodule












































 // FUNCTIONAL































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_POWER_LVC_WPAD_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_refgen: The REFGEN block (sky130_fd_io__top_refgen) is used to
 *             provide the input trip point (VINREF) for the
 *             differential input buffer in SIO and also
 *             the output buffer regulated output level (VOUTREF).
 *             Verilog HDL for "sky130_fd_io",
 *             "sky130_fd_io_top_refgen" "behavioral_tmp".
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_refgen (VINREF, VOUTREF, REFLEAK_BIAS,
                                 VCCD, VCCHIB, VDDA, VDDIO, VDDIO_Q, VSSD, VSSIO, VSSIO_Q,
                                 HLD_H_N, IBUF_SEL, OD_H, VOHREF, VREF_SEL, VREG_EN, VTRIP_SEL);
wire error_vsel;
output VINREF;
output VOUTREF;
inout REFLEAK_BIAS;
inout VCCD;
inout VCCHIB;
inout VDDA;
inout VDDIO;
inout VDDIO_Q;
inout VSSD;
inout VSSIO;
inout VSSIO_Q;
input HLD_H_N;
input IBUF_SEL;
input OD_H;
input VOHREF;
input VREF_SEL;
input VREG_EN;
input VTRIP_SEL;
reg [2:0] dm_final;
reg       slow_final, vtrip_sel_final, inp_dis_final, hld_ovr_final;
reg [2:0] dm;
reg       slow, inp_dis, hld_ovr;
reg [1:0] vsel;
wire  pwr_good_active_mode    = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0)    && (VCCD===1);
wire  pwr_good_hold_mode      = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0);
always @(*)
begin
    if (^OD_H===1'bx || !pwr_good_hold_mode || (OD_H===0 && ^HLD_H_N===1'bx))
    begin
        dm_final 	= 3'bxxx;
        slow_final 	= 1'bx;
        vtrip_sel_final	= 1'bx;
        inp_dis_final 	= 1'bx;
        hld_ovr_final 	= 1'bx;
    end
    else if (OD_H===1)
    begin
        dm_final 	= 3'b000;
        slow_final 	= 1'b0;
        vtrip_sel_final	= 1'b0;
        inp_dis_final 	= 1'b0;
        hld_ovr_final 	= 1'b0;
    end
    else if (HLD_H_N===1)
    begin
        dm_final 	= (^dm[2:0] === 1'bx	|| !pwr_good_active_mode) ? 3'bxxx : dm;
        slow_final 	= (^slow 	=== 1'bx	|| !pwr_good_active_mode) ? 1'bx   : slow;
        vtrip_sel_final	= (^VTRIP_SEL 	=== 1'bx	|| !pwr_good_active_mode) ? 1'bx   : VTRIP_SEL;
        inp_dis_final 	= (^inp_dis	=== 1'bx	|| !pwr_good_active_mode) ? 1'bx   : inp_dis;
        hld_ovr_final 	= (^hld_ovr 	=== 1'bx	|| !pwr_good_active_mode) ? 1'bx   : hld_ovr;
    end
end
reg dis_err_msgs;
initial
begin
    dis_err_msgs = 1'b1;


    #1;
    dis_err_msgs = 1'b0;

end
assign error_vsel = (vsel[1]===1 && vsel[0]===1);
always @(*)
begin
    if (!dis_err_msgs)
    begin
        if (error_vsel==1) $display(" ===ERROR=== sky130_fd_io__top_refgen : %m : Incorrect inputs on vsel[1:0] = 11",$stime);
    end
end
endmodule






























































































 // FUNCTIONAL































































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_REFGEN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_refgen_new: The REFGEN block (sky130_fd_io__top_refgen) is used
 *                 to provide the input trip point (VINREF) for the
 *                 differential input buffer in SIO and also
 *                 the output buffer regulated output level (VOUTREF).
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_refgen_new (VINREF, VOUTREF, REFLEAK_BIAS,
                                     VCCD, VCCHIB, VDDA, VDDIO, VDDIO_Q, VSSD, VSSIO, VSSIO_Q, VSWITCH, VSSA,
                                     AMUXBUS_A, AMUXBUS_B, DFT_REFGEN, HLD_H_N, IBUF_SEL, ENABLE_H, ENABLE_VDDA_H, VOH_SEL, VOHREF,
                                     VREF_SEL, VREG_EN, VTRIP_SEL, VOUTREF_DFT, VINREF_DFT);
output VINREF;
output VOUTREF;
inout REFLEAK_BIAS;
inout VCCD;
inout VCCHIB;
inout VDDA;
inout VDDIO;
inout VDDIO_Q;
inout VSSD;
inout VSSIO;
inout VSSIO_Q;
inout VSWITCH;
inout VSSA;
inout AMUXBUS_A;
inout AMUXBUS_B;
input DFT_REFGEN;
input HLD_H_N;
input IBUF_SEL;
input ENABLE_H;
input ENABLE_VDDA_H;
input [2:0] VOH_SEL;
input VOHREF;
input [1:0] VREF_SEL;
input VREG_EN;
input VTRIP_SEL;
inout VOUTREF_DFT;
inout VINREF_DFT;
reg ibuf_sel_final, vtrip_sel_final, vreg_en_final, dft_refgen_final, vref_sel_int_final;
reg [2:0] voh_sel_final;
reg [1:0] vref_sel_final;
reg vohref_int;
wire  pwr_good_active_mode_1    = (VDDIO_Q===1) && (VSSD===0) && (VCCD===1);
wire  pwr_good_hold_mode_1      = (VDDIO_Q===1) && (VSSD===0);
wire  pwr_good_hold_mode_2   	= (VDDA===1) && (VSWITCH===1) && (VSSA===0) && (VSSD===0);
wire  pwr_good_active_mode_2 	= (VDDA===1) && (VSWITCH===1) && (VSSA===0) && (VSSD===0) && (VCCD===1);
wire  pwr_good_hold_mode_3   	= (VSWITCH===1) && (VSSD===0) && (VSSA===0);
wire  pwr_good_active_mode_3 	= (VSWITCH===1) && (VSSD===0) && (VCCD===1) && (VSSA===0);




parameter STARTUP_TIME_VOUTREF = 50000;
parameter STARTUP_TIME_VINREF  = 50000;

integer startup_time_vinref,startup_time_voutref;
initial begin
    startup_time_vinref 	= vref_sel_int_final===1 && vtrip_sel_final===0 ? STARTUP_TIME_VINREF : 0;
    startup_time_voutref 	= STARTUP_TIME_VOUTREF;
end
wire 	notifier_enable_h, notifier_vtrip_sel, notifier_ibuf_sel, notifier_vref_sel,
      notifier_voh_sel, notifier_vreg_en, notifier_dft_refgen, notifier_vref_sel_int;
always @(*)
begin : LATCH_ibuf_sel
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode_1 || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        ibuf_sel_final 		<= 1'bx;
    else if (ENABLE_H===0)
        ibuf_sel_final 		<= 1'b0;
    else if (HLD_H_N===1)
        ibuf_sel_final 		<= (^IBUF_SEL 	  === 1'bx  || !pwr_good_active_mode_1) ? 1'bx 	: IBUF_SEL;
end
always @(notifier_enable_h or notifier_ibuf_sel)
begin
    disable LATCH_ibuf_sel; ibuf_sel_final <= 1'bx;
end
always @(*)
begin : LATCH_vtrip_sel
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode_1 || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        vtrip_sel_final 		<= 1'bx;
    else if (ENABLE_H===0)
        vtrip_sel_final 		<= 1'b0;
    else if (HLD_H_N===1)
        vtrip_sel_final 		<= (^VTRIP_SEL 	  === 1'bx  || !pwr_good_active_mode_1) ? 1'bx 	: VTRIP_SEL;
end
always @(notifier_enable_h or notifier_vtrip_sel)
begin
    disable LATCH_vtrip_sel; vtrip_sel_final <= 1'bx;
end
always @(*)
begin : LATCH_vreg_en
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode_1 || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        vreg_en_final 		<= 1'bx;
    else if (ENABLE_H===0)
        vreg_en_final 		<= 1'b0;
    else if (HLD_H_N===1)
        vreg_en_final 		<= (^VREG_EN 	  === 1'bx  || !pwr_good_active_mode_1) ? 1'bx 	: VREG_EN;
end
always @(notifier_enable_h or notifier_vreg_en)
begin
    disable LATCH_vreg_en; vreg_en_final <= 1'bx;
end
always @(*)
begin : LATCH_vref_sel_int
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode_1 || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        vref_sel_int_final 		<= 1'bx;
    else if (ENABLE_H===0)
        vref_sel_int_final 		<= 1'b0;
    else if (HLD_H_N===1)
        vref_sel_int_final 		<= (^VREF_SEL[1:0]  === 1'bx  || !pwr_good_active_mode_1) ? 1'bx : (VREF_SEL[1] || VREF_SEL[0]);
end
always @(notifier_enable_h or notifier_vref_sel_int)
begin
    disable LATCH_vref_sel; vref_sel_int_final <= 1'bx;
end
always @(*)
begin : LATCH_vref_sel
    if (^ENABLE_VDDA_H===1'bx || ^ENABLE_H===1'bx ||!pwr_good_hold_mode_2 || (ENABLE_VDDA_H===1 && ENABLE_H===1 && ^HLD_H_N===1'bx))
        vref_sel_final 	= 2'bxx;
    else if (ENABLE_VDDA_H===0 || ENABLE_H===0)
        vref_sel_final	= 2'b00;
    else if (HLD_H_N===1)
        vref_sel_final 	= (^VREF_SEL[1:0]=== 1'bx || !pwr_good_active_mode_2) ? 2'bxx : VREF_SEL;
end
always @(notifier_enable_h or notifier_vref_sel)
begin
    disable LATCH_vref_sel; vref_sel_final <= 2'bxx;
end
always @(*)
begin : LATCH_dft_refgen
    if (^ENABLE_VDDA_H===1'bx || ^ENABLE_H===1'bx ||!pwr_good_hold_mode_2 || (ENABLE_VDDA_H===1 && ENABLE_H===1 &&^HLD_H_N===1'bx))
        dft_refgen_final 	= 2'bxx;
    else if (ENABLE_VDDA_H===0 || ENABLE_H===0)
        dft_refgen_final	= 2'b00;
    else if (HLD_H_N===1)
        dft_refgen_final 	= (^DFT_REFGEN=== 1'bx || !pwr_good_active_mode_2) ? 2'bxx : DFT_REFGEN;
end
always @(notifier_enable_h or notifier_dft_refgen)
begin
    disable LATCH_dft_refgen; dft_refgen_final <= 2'bxx;
end
always @(*)
begin : LATCH_voh_sel
    if (^ENABLE_VDDA_H===1'bx ||^ENABLE_H===1'bx || !pwr_good_hold_mode_3 || (ENABLE_VDDA_H===1 && ENABLE_H===1 && ^HLD_H_N===1'bx))
        voh_sel_final 	= 3'bxxx;
    else if (ENABLE_VDDA_H===0 || ENABLE_H===0)
        voh_sel_final	= 3'b000;
    else if (HLD_H_N===1)
        voh_sel_final 	= (^VOH_SEL[2:0]=== 1'bx || !pwr_good_active_mode_3) ? 3'bxxx : VOH_SEL;
end
always @(notifier_enable_h or notifier_voh_sel)
begin
    disable LATCH_voh_sel; voh_sel_final <= 2'bxx;
end
always @(*)
begin
    case (vref_sel_final[1:0])
        2'b00, 2'b01   : vohref_int = VOHREF!==1'b1 ? 1'bx : VOHREF;
        2'b10	       : vohref_int = ^AMUXBUS_A!==1'b1 ? 1'bx : AMUXBUS_A;
        2'b11	       : vohref_int = ^AMUXBUS_B!==1'b1 ? 1'bx : AMUXBUS_B;
        default	       : vohref_int = 1'bx;
    endcase
end
wire vohref_final = ENABLE_VDDA_H===1'b1 ? vohref_int : 1'bx;
assign #(startup_time_voutref,0) VOUTREF = (REFLEAK_BIAS===1'bx) ? 1'bx : (REFLEAK_BIAS===1 ? vohref_final:1'bz);
assign VOUTREF_DFT = dft_refgen_final===1 ? VOUTREF : (dft_refgen_final===0 ? 1'bz : 1'bx);
assign REFLEAK_BIAS = VCCHIB!==1 ? 1'bx : (vreg_en_final || (ibuf_sel_final && vref_sel_int_final));
reg vinref_tmp;
always @(*)
begin
    if (ibuf_sel_final===1'bx
            || (ibuf_sel_final===1 && (vref_sel_int_final===1'bx || vtrip_sel_final===1'bx))
            || (ibuf_sel_final===1 && vref_sel_int_final===1 && (VCCHIB!==1 || vohref_int!==1))
            || (ibuf_sel_final===1 && vref_sel_int_final===1 && vtrip_sel_final===0 && ^voh_sel_final[2:0]===1'bx))
        vinref_tmp = 1'bx;
    else
        vinref_tmp = ibuf_sel_final===0 ? 1'bz : 1'b1;
end
assign #(startup_time_vinref,0) VINREF = vinref_tmp;
assign VINREF_DFT = dft_refgen_final===1 ? VINREF : (dft_refgen_final===0 ? 1'bz : 1'bx);
endmodule
































































































































































































 // FUNCTIONAL



































































































































































































































































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_REFGEN_NEW_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_sio: Special I/O PAD that provides additionally a
 *          regulated output buffer and a differential input buffer.
 *          SIO cells are ONLY available IN pairs (see top_sio_macro).
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_sio (IN_H, PAD_A_NOESD_H, PAD, DM, HLD_H_N, INP_DIS, IN,
                              ENABLE_H, OE_N, SLOW, VTRIP_SEL, VINREF, VOUTREF, VREG_EN, IBUF_SEL,
                              REFLEAK_BIAS, PAD_A_ESD_0_H, TIE_LO_ESD, HLD_OVR, OUT,
                              PAD_A_ESD_1_H
                              ,VSSIO, VSSIO_Q, VSSD, VCCD, VDDIO, VCCHIB, VDDIO_Q
                             );
output IN_H;
inout PAD_A_NOESD_H;
inout PAD;
input [2:0] DM;
input HLD_H_N;
input INP_DIS;
output IN;
input ENABLE_H;
input OE_N;
input SLOW;
input VTRIP_SEL;
input VINREF;
input VOUTREF;
input VREG_EN;
input IBUF_SEL;
input REFLEAK_BIAS;
inout PAD_A_ESD_0_H;
output TIE_LO_ESD;
input HLD_OVR;
input OUT;
inout PAD_A_ESD_1_H;
inout VSSIO;
inout VSSIO_Q;
inout VSSD;
inout VCCD;
inout VDDIO;
inout VCCHIB;
inout VDDIO_Q;
reg [2:0] dm_final;
reg slow_final, vtrip_sel_final, inp_dis_final, out_final, oe_n_final, hld_ovr_final;
reg ibuf_sel_final, vreg_en_final;
wire notifier_dm, notifier_slow, notifier_oe_n, notifier_out, notifier_vtrip_sel, notifier_hld_ovr, notifier_inp_dis, notifier_vreg_en,notifier_ibuf_sel;
wire notifier_enable_h;
wire  pwr_good_hold_ovr_mode  = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0)    && (VCCHIB===1);
wire  pwr_good_active_mode    = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0)    && (VCCD===1);
wire  pwr_good_hold_mode      = (VDDIO_Q===1) && (VDDIO===1)  && (VSSD===0);
wire  pwr_good_inpbuff_lv     = (VDDIO_Q===1) && (VCCHIB===1) && (VSSD===0)    && (VDDIO===1) && (VSSIO===0);
wire  pwr_good_inpbuff_hv     = (VDDIO_Q===1) && (VSSD===0)   && (VDDIO===1) && (VSSIO===0);
wire  pwr_good_output_driver  = (VDDIO===1)   && (VDDIO_Q===1)&& (VSSIO===0)   && (VSSD===0);
wire pad_tristate = oe_n_final === 1 || dm_final === 3'b000 || dm_final === 3'b001;
wire x_on_pad  =  !pwr_good_output_driver
     || (dm_final !== 3'b000 && dm_final !== 3'b001 && oe_n_final===1'bx)
     || (^dm_final[2:0] === 1'bx && oe_n_final===1'b0)
     || (slow_final===1'bx && dm_final !== 3'b000 && dm_final !== 3'b001 && oe_n_final===1'b0)
     || (vreg_en_final===1'bx && dm_final !== 3'b000 && dm_final !== 3'b001 && oe_n_final===1'b0)
     || ((VOUTREF!==1'b1 || REFLEAK_BIAS!==1'b1) && vreg_en_final===1'b1 && dm_final !== 3'b000 && dm_final !== 3'b001 && oe_n_final===1'b0 );




parameter SLOW_1_DELAY= 0;
parameter SLOW_0_DELAY= 0;

integer slow_1_delay,slow_0_delay,slow_delay;
initial slow_1_delay = SLOW_1_DELAY;
initial slow_0_delay = SLOW_0_DELAY;
always @(*)
begin
    if (SLOW===1)
        slow_delay = slow_1_delay;
    else
        slow_delay = slow_0_delay;
end
bufif1 (pull1, strong0) #slow_delay  dm2 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b010));
bufif1 (strong1, pull0)  #slow_delay dm3 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b011));
bufif1 (highz1, strong0) #slow_delay dm4 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b100));
bufif1 (strong1, highz0) #slow_delay dm5 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b101));
bufif1 (strong1, strong0)#slow_delay dm6 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b110));
bufif1 (pull1, pull0)   #slow_delay  dm7 (PAD, out_final, x_on_pad===1 ? 1'bx : (pad_tristate===0 && dm_final===3'b111));
tran pad_esd_1 (PAD,PAD_A_NOESD_H);
tran pad_esd_2 (PAD,PAD_A_ESD_0_H);
tran pad_esd_3 (PAD,PAD_A_ESD_1_H);
wire x_on_in  =  (pwr_good_inpbuff_hv===0)
     || (inp_dis_final===1'bx    && dm_final !== 3'b000)
     || (inp_dis_final===0 	     && ^dm_final[2:0] === 1'bx )
     || (vtrip_sel_final===1'bx  && inp_dis_final===0  && dm_final !== 3'b000)
     || (ibuf_sel_final===1'bx   && inp_dis_final===0  && dm_final !== 3'b000)
     || (VINREF!==1'b1  && inp_dis_final===0  && dm_final !== 3'b000 && ibuf_sel_final===1);
wire disable_inp_buff = (dm_final===3'b000 || inp_dis_final===1);
assign IN_H = x_on_in===1 ? 1'bx : (disable_inp_buff===1 ? 0 : (^PAD===1'bx ? 1'bx : PAD));
assign IN = pwr_good_inpbuff_lv===1 ? IN_H : 1'bx;
assign TIE_LO_ESD = VSSIO===1'b0 ? 1'b0 : 1'bx;
always @(*)
begin : LATCH_dm
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        dm_final 	<= 3'bxxx;
    else if (ENABLE_H===0)
        dm_final 	<= 3'b000;
    else if (HLD_H_N===1)
        dm_final 	<= (^DM[2:0]	=== 1'bx	|| !pwr_good_active_mode) ? 3'bxxx : DM;
end
always @(notifier_enable_h or notifier_dm)
begin
    disable LATCH_dm; dm_final <= 3'bxxx;
end
always @(*)
begin : LATCH_inp_dis
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        inp_dis_final 	<= 1'bx;
    else if (ENABLE_H===0)
        inp_dis_final 	<= 1'b0;
    else if (HLD_H_N===1)
        inp_dis_final 	<= (^INP_DIS === 1'bx	|| !pwr_good_active_mode) ? 1'bx : INP_DIS;
end
always @(notifier_enable_h or notifier_inp_dis)
begin
    disable LATCH_inp_dis; inp_dis_final <= 1'bx;
end
always @(*)
begin : LATCH_vtrip_sel
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        vtrip_sel_final 	<= 1'bx;
    else if (ENABLE_H===0)
        vtrip_sel_final 	<= 1'b0;
    else if (HLD_H_N===1)
        vtrip_sel_final 	<= (^VTRIP_SEL === 1'bx	|| !pwr_good_active_mode) ? 1'bx : VTRIP_SEL;
end
always @(notifier_enable_h or notifier_vtrip_sel)
begin
    disable LATCH_vtrip_sel; vtrip_sel_final <= 1'bx;
end
always @(*)
begin : LATCH_slow
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        slow_final 	<= 1'bx;
    else if (ENABLE_H===0)
        slow_final 	<= 1'b0;
    else if (HLD_H_N===1)
        slow_final 	<= (^SLOW === 1'bx	|| !pwr_good_active_mode) ? 1'bx : SLOW;
end
always @(notifier_enable_h or notifier_slow)
begin
    disable LATCH_slow; slow_final <= 1'bx;
end
always @(*)
begin : LATCH_hld_ovr
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        hld_ovr_final 	<= 1'bx;
    else if (ENABLE_H===0)
        hld_ovr_final 	<= 1'b0;
    else if (HLD_H_N===1)
        hld_ovr_final 	<= (^HLD_OVR === 1'bx	|| !pwr_good_active_mode) ? 1'bx : HLD_OVR;
end
always @(notifier_enable_h or notifier_hld_ovr)
begin
    disable LATCH_hld_ovr; hld_ovr_final <= 1'bx;
end
always @(*)
begin : LATCH_vreg_en
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        vreg_en_final 	<= 1'bx;
    else if (ENABLE_H===0)
        vreg_en_final 	<= 1'b0;
    else if (HLD_H_N===1)
        vreg_en_final 	<= (^VREG_EN === 1'bx	|| !pwr_good_active_mode) ? 1'bx : VREG_EN;
end
always @(notifier_enable_h or notifier_vreg_en)
begin
    disable LATCH_vreg_en; vreg_en_final <= 1'bx;
end
always @(*)
begin : LATCH_ibuf_sel
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && ^HLD_H_N===1'bx))
        ibuf_sel_final 	<= 1'bx;
    else if (ENABLE_H===0)
        ibuf_sel_final 	<= 1'b0;
    else if (HLD_H_N===1)
        ibuf_sel_final 	<= (^IBUF_SEL === 1'bx	|| !pwr_good_active_mode) ? 1'bx : IBUF_SEL;
end
always @(notifier_enable_h or notifier_ibuf_sel)
begin
    disable LATCH_ibuf_sel; ibuf_sel_final <= 1'bx;
end
always @(*)
begin : LATCH_oe_n
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && (^HLD_H_N===1'bx || (HLD_H_N===0 && hld_ovr_final===1'bx))))
        oe_n_final 	<= 1'bx;
    else if (ENABLE_H===0)
        oe_n_final 	<= 1'b0;
    else if (HLD_H_N===1 || hld_ovr_final===1)
        oe_n_final  	<= (^OE_N  === 1'bx  || !pwr_good_hold_ovr_mode) ? 1'bx   : OE_N;
end
always @(notifier_enable_h or notifier_oe_n)
begin
    disable LATCH_oe_n; oe_n_final <= 1'bx;
end
always @(*)
begin : LATCH_out
    if (^ENABLE_H===1'bx || !pwr_good_hold_mode || (ENABLE_H===1 && (^HLD_H_N===1'bx || (HLD_H_N===0 && hld_ovr_final===1'bx))))
        out_final 	<= 1'bx;
    else if (ENABLE_H===0)
        out_final 	<= 1'b0;
    else if (HLD_H_N===1 || hld_ovr_final===1)
        out_final  	<= (^OUT  === 1'bx  || !pwr_good_hold_ovr_mode) ? 1'bx   : OUT;
end
always @(notifier_enable_h or notifier_out)
begin
    disable LATCH_out; out_final <= 1'bx;
end
reg dis_err_msgs;
initial
begin
    dis_err_msgs = 1'b1;


    #1;
    dis_err_msgs = 1'b0;

end
always @(*)
begin
    if (!dis_err_msgs)
    begin
        if (vreg_en_final===1 && (dm_final!==3'b011 && dm_final!==3'b110 && dm_final!==3'b101))
            $display(" ===INFO=== sky130_fd_io__top_sio :  In regulated output driver mode (vreg_en_final=1), dm_final should be either \011 / 101 / 110 (i.E.strong-pullup mode) inorder for regulated mode to be effective : DM (= %b) and VREG_EN (= %b): %m",dm_final,vreg_en_final,$stime);
    end
end
endmodule



















































































































































































































































 // FUNCTIONAL









































































































































































































































































































































































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_SIO_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_sio_macro: sky130_fd_io__sio_macro consists of two SIO cells
 *                and a reference generator cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_sio_macro (
           VCCD,
           VCCHIB,
           VDDA,
           VDDIO,
           VDDIO_Q,
           VSSD,
           VSSIO,
           VSSIO_Q,
           VSWITCH,
           VSSA,
           IN,
           IN_H,
           TIE_LO_ESD,
           AMUXBUS_A,
           AMUXBUS_B,
           PAD,
           PAD_A_ESD_0_H,
           PAD_A_ESD_1_H,
           PAD_A_NOESD_H,
           VINREF_DFT,
           VOUTREF_DFT,
           DFT_REFGEN,
           DM0,
           DM1,
           HLD_H_N,
           HLD_H_N_REFGEN,
           HLD_OVR,
           IBUF_SEL,
           IBUF_SEL_REFGEN,
           INP_DIS,
           ENABLE_H,
           ENABLE_VDDA_H,
           OE_N,
           OUT,
           SLOW,
           VOH_SEL,
           VOHREF,
           VREF_SEL,
           VREG_EN,
           VREG_EN_REFGEN,
           VTRIP_SEL,
           VTRIP_SEL_REFGEN
       );
wire VOUTREF;
wire VINREF;
wire REFLEAK_BIAS;
inout VCCD;
inout VCCHIB;
inout VDDA;
inout VDDIO;
inout VDDIO_Q;
inout VSSD;
inout VSSIO;
inout VSSIO_Q;
inout VSWITCH;
inout VSSA;
inout AMUXBUS_A;
inout AMUXBUS_B;
inout VINREF_DFT;
inout VOUTREF_DFT;
input DFT_REFGEN;
input HLD_H_N_REFGEN;
input IBUF_SEL_REFGEN;
input ENABLE_VDDA_H;
input ENABLE_H;
input VOHREF;
input VREG_EN_REFGEN;
input VTRIP_SEL_REFGEN;
output [1:0]  TIE_LO_ESD;
output [1:0]  IN_H;
output [1:0]  IN;
inout [1:0]  PAD_A_NOESD_H;
inout [1:0]  PAD;
inout [1:0]  PAD_A_ESD_1_H;
inout [1:0]  PAD_A_ESD_0_H;
input [1:0]  SLOW;
input [1:0]  VTRIP_SEL;
input [1:0]  HLD_H_N;
input [1:0]  VREG_EN;
input [2:0]  VOH_SEL;
input [1:0]  INP_DIS;
input [1:0]  HLD_OVR;
input [1:0]  OE_N;
input [1:0]  VREF_SEL;
input [1:0]  IBUF_SEL;
input [2:0]  DM0;
input [2:0]  DM1;
input [1:0]  OUT;
reg 	notifier_enable_h_refgen,
     notifier_vtrip_sel_refgen,
     notifier_vreg_en_refgen,
     notifier_ibuf_sel_refgen,
     notifier_vref_sel,
     notifier_vref_sel_int,
     notifier_voh_sel,
     notifier_dft_refgen;
reg	 notifier_enable_h_0;
reg	 notifier_hld_ovr_0;
reg	 notifier_dm_0;
reg	 notifier_inp_dis_0;
reg	 notifier_vtrip_sel_0;
reg	 notifier_slow_0;
reg	 notifier_oe_n_0;
reg	 notifier_out_0;
reg	 notifier_vreg_en_0;
reg	 notifier_ibuf_sel_0;
reg	 notifier_enable_h_1;
reg	 notifier_hld_ovr_1;
reg	 notifier_dm_1;
reg	 notifier_inp_dis_1;
reg	 notifier_vtrip_sel_1;
reg	 notifier_slow_1;
reg	 notifier_oe_n_1;
reg	 notifier_out_1;
reg	 notifier_vreg_en_1;
reg	 notifier_ibuf_sel_1;
wire enable_vdda_h_and_enable_h = ENABLE_VDDA_H==1'b1 && ENABLE_H==1'b1;
sky130_fd_io__top_refgen_new REFGEN (
                                 .VSWITCH                                      (VSWITCH),
                                 .VSSIO_Q                                      (VSSIO_Q),
                                 .VDDIO_Q                                      (VDDIO_Q),
                                 .VSSIO                                        (VSSIO),
                                 .VSSD                                         (VSSD),
                                 .VCCHIB                                       (VCCHIB),
                                 .VDDIO                                        (VDDIO),
                                 .VCCD                                         (VCCD),
                                 .VDDA                                         (VDDA),
                                 .VSSA					  (VSSA),
                                 .VOH_SEL                                      (VOH_SEL[2:0]),
                                 .VREF_SEL                                     (VREF_SEL[1:0]),
                                 .VOHREF                                       (VOHREF),
                                 .VINREF_DFT                                   (VINREF_DFT),
                                 .VOUTREF_DFT                                  (VOUTREF_DFT),
                                 .DFT_REFGEN                                   (DFT_REFGEN),
                                 .AMUXBUS_A                                    (AMUXBUS_A),
                                 .AMUXBUS_B                                    (AMUXBUS_B),
                                 .VOUTREF                                      (VOUTREF),
                                 .VREG_EN                                      (VREG_EN_REFGEN),
                                 .IBUF_SEL                                     (IBUF_SEL_REFGEN),
                                 .VINREF                                       (VINREF),
                                 .VTRIP_SEL                                    (VTRIP_SEL_REFGEN),
                                 .ENABLE_H					  (ENABLE_H),
                                 .ENABLE_VDDA_H				  (ENABLE_VDDA_H),
                                 .HLD_H_N                                      (HLD_H_N_REFGEN),
                                 .REFLEAK_BIAS                                 (REFLEAK_BIAS)
                             );
sky130_fd_io__top_sio SIO_PAIR_1_ (
                          .VDDIO                                        (VDDIO),
                          .VCCD                                         (VCCD),
                          .VDDIO_Q                                      (VDDIO_Q),
                          .VCCHIB                                       (VCCHIB),
                          .VSSIO                                        (VSSIO),
                          .VSSIO_Q                                      (VSSIO_Q),
                          .VSSD                                         (VSSD),
                          .PAD                                          (PAD[1]),
                          .IN_H                                         (IN_H[1]),
                          .DM                                           (DM1[2:0]),
                          .HLD_H_N                                      (HLD_H_N[1]),
                          .PAD_A_ESD_1_H                                (PAD_A_ESD_1_H[1]),
                          .PAD_A_ESD_0_H                                (PAD_A_ESD_0_H[1]),
                          .ENABLE_H                                     (ENABLE_H),
                          .OUT                                          (OUT[1]),
                          .OE_N                                         (OE_N[1]),
                          .SLOW                                         (SLOW[1]),
                          .VTRIP_SEL                                    (VTRIP_SEL[1]),
                          .INP_DIS                                      (INP_DIS[1]),
                          .TIE_LO_ESD                                   (TIE_LO_ESD[1]),
                          .IN                                           (IN[1]),
                          .VINREF                                       (VINREF),
                          .VOUTREF                                      (VOUTREF),
                          .REFLEAK_BIAS                                 (REFLEAK_BIAS),
                          .PAD_A_NOESD_H                                (PAD_A_NOESD_H[1]),
                          .VREG_EN                                      (VREG_EN[1]),
                          .IBUF_SEL                                     (IBUF_SEL[1]),
                          .HLD_OVR                                      (HLD_OVR[1])
                      );
sky130_fd_io__top_sio SIO_PAIR_0_ (
                          .VDDIO                                        (VDDIO),
                          .VCCD                                         (VCCD),
                          .VDDIO_Q                                      (VDDIO_Q),
                          .VCCHIB                                       (VCCHIB),
                          .VSSIO                                        (VSSIO),
                          .VSSIO_Q                                      (VSSIO_Q),
                          .VSSD                                         (VSSD),
                          .PAD                                          (PAD[0]),
                          .IN_H                                         (IN_H[0]),
                          .DM                                           (DM0[2:0]),
                          .HLD_H_N                                      (HLD_H_N[0]),
                          .PAD_A_ESD_1_H                                (PAD_A_ESD_1_H[0]),
                          .PAD_A_ESD_0_H                                (PAD_A_ESD_0_H[0]),
                          .ENABLE_H                                     (ENABLE_H),
                          .OUT                                          (OUT[0]),
                          .OE_N                                         (OE_N[0]),
                          .SLOW                                         (SLOW[0]),
                          .VTRIP_SEL                                    (VTRIP_SEL[0]),
                          .INP_DIS                                      (INP_DIS[0]),
                          .TIE_LO_ESD                                   (TIE_LO_ESD[0]),
                          .IN                                           (IN[0]),
                          .VINREF                                       (VINREF),
                          .VOUTREF                                      (VOUTREF),
                          .REFLEAK_BIAS                                 (REFLEAK_BIAS),
                          .PAD_A_NOESD_H                                (PAD_A_NOESD_H[0]),
                          .VREG_EN                                      (VREG_EN[0]),
                          .IBUF_SEL                                     (IBUF_SEL[0]),
                          .HLD_OVR                                      (HLD_OVR[0])
                      );
endmodule





























































































































































































































































































































































































































































































 // FUNCTIONAL

































































































































































































































































































































































































































































































































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_SIO_MACRO_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * top_xres4v2: XRES (Input buffer with Glitch filter).
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_fd_io__top_xres4v2 ( TIE_WEAK_HI_H,  XRES_H_N, TIE_HI_ESD, TIE_LO_ESD,
                                   AMUXBUS_A, AMUXBUS_B, PAD, PAD_A_ESD_H, ENABLE_H, EN_VDDIO_SIG_H, INP_SEL_H, FILT_IN_H,
                                   DISABLE_PULLUP_H, PULLUP_H, ENABLE_VDDIO
                                   ,VCCD, VCCHIB, VDDA, VDDIO,VDDIO_Q, VSSA, VSSD, VSSIO, VSSIO_Q, VSWITCH
                                 );
output XRES_H_N;
inout AMUXBUS_A;
inout AMUXBUS_B;
inout PAD;
input DISABLE_PULLUP_H;
input ENABLE_H;
input EN_VDDIO_SIG_H;
input INP_SEL_H;
input FILT_IN_H;
inout PULLUP_H;
input ENABLE_VDDIO;
input VCCD;
input VCCHIB;
input VDDA;
input VDDIO;
input VDDIO_Q;
input VSSA;
input VSSD;
input VSSIO;
input VSSIO_Q;
input VSWITCH;
wire mode_vcchib;
wire pwr_good_xres_tmp 	= (VDDIO===1) && (VDDIO_Q===1) && ((mode_vcchib && ENABLE_VDDIO)===1 ? VCCHIB===1 : 1'b1) &&  (VSSIO===0) && (VSSD===0);
wire pwr_good_xres_h_n 		= (VDDIO_Q===1) && (VSSD===0);
wire pwr_good_pullup 		= (VDDIO===1) && (VSSD===0);
inout PAD_A_ESD_H;
output TIE_HI_ESD;
output TIE_LO_ESD;
inout TIE_WEAK_HI_H;
wire tmp1;
pullup (pull1) p1 (tmp1); tranif1 x_pull_1 (TIE_WEAK_HI_H, tmp1, pwr_good_pullup===0  ? 1'bx : 1);
tran p2 (PAD, PAD_A_ESD_H);
buf p4 (TIE_HI_ESD, VDDIO);
buf p5 (TIE_LO_ESD, VSSIO);
wire tmp;
pullup (pull1) p3 (tmp); tranif0 x_pull (PULLUP_H, tmp, pwr_good_pullup===0 || ^DISABLE_PULLUP_H===1'bx ? 1'bx : DISABLE_PULLUP_H);
parameter MAX_WARNING_COUNT = 100;




parameter MIN_DELAY = 50;
parameter MAX_DELAY = 600;

integer min_delay, max_delay;
initial begin
    min_delay = MIN_DELAY;
    max_delay = MAX_DELAY;
end



parameter DISABLE_ENABLE_VDDIO_CHANGE_X = 0;

integer     disable_enable_vddio_change_x    = DISABLE_ENABLE_VDDIO_CHANGE_X;
reg notifier_enable_h;
specify



    specparam DELAY = 50;

    if (INP_SEL_H==0  &  ENABLE_H==0  & ENABLE_VDDIO==0 & EN_VDDIO_SIG_H==1) (PAD   => XRES_H_N) =  (0:0:0 , 0:0:0);
    if (INP_SEL_H==0  &  ENABLE_H==1  & ENABLE_VDDIO==1 & EN_VDDIO_SIG_H==1) (PAD   => XRES_H_N) =  (0:0:0 , 0:0:0);
    if (INP_SEL_H==0  &  ENABLE_H==1  & ENABLE_VDDIO==1 & EN_VDDIO_SIG_H==0) (PAD   => XRES_H_N) =  (0:0:0 , 0:0:0);
    if (INP_SEL_H==0  &  ENABLE_H==0  & ENABLE_VDDIO==0 & EN_VDDIO_SIG_H==0) (PAD   => XRES_H_N) =  (0:0:0 , 0:0:0);
    if (INP_SEL_H==1) (FILT_IN_H => XRES_H_N) =  (0:0:0 , 0:0:0);
    specparam tsetup = 0;
    specparam thold = 5;
endspecify
reg corrupt_enable;
always @(notifier_enable_h)
begin
    corrupt_enable <= 1'bx;
end
initial
begin
    corrupt_enable = 1'b0;
end
always @(PAD or ENABLE_H or EN_VDDIO_SIG_H or ENABLE_VDDIO or INP_SEL_H or FILT_IN_H or pwr_good_xres_tmp or DISABLE_PULLUP_H or PULLUP_H or TIE_WEAK_HI_H)
begin
    corrupt_enable <= 1'b0;
end
assign mode_vcchib 	= ENABLE_H && !EN_VDDIO_SIG_H;
wire xres_tmp 	= (pwr_good_xres_tmp===0 || ^PAD===1'bx || (mode_vcchib===1'bx ) ||(mode_vcchib!==1'b0 && ^ENABLE_VDDIO===1'bx) || (corrupt_enable===1'bx) ||
                  (mode_vcchib===1'b1 && ENABLE_VDDIO===0 && (disable_enable_vddio_change_x===0)))
     ? 1'bx : PAD;
wire x_on_xres_h_n = (pwr_good_xres_h_n===0
                      || ^INP_SEL_H===1'bx
                      || INP_SEL_H===1 && ^FILT_IN_H===1'bx
                      || INP_SEL_H===0 && xres_tmp===1'bx);
assign #1  XRES_H_N = x_on_xres_h_n===1 ? 1'bx : (INP_SEL_H===1 ? FILT_IN_H : xres_tmp);
realtime t_pad_current_transition,t_pad_prev_transition;
realtime t_filt_in_h_current_transition,t_filt_in_h_prev_transition;
realtime pad_pulse_width, filt_in_h_pulse_width;
always @(PAD)
begin
    if (^PAD !== 1'bx)
    begin
        t_pad_prev_transition    	= t_pad_current_transition;
        t_pad_current_transition 	= $realtime;
        pad_pulse_width 	     	= t_pad_current_transition - t_pad_prev_transition;
    end
    else
    begin
        t_pad_prev_transition 		= 0;
        t_pad_current_transition 	= 0;
        pad_pulse_width 		= 0;
    end
end
always @(FILT_IN_H)
begin
    if (^FILT_IN_H !== 1'bx)
    begin
        t_filt_in_h_prev_transition    			= t_filt_in_h_current_transition;
        t_filt_in_h_current_transition 			= $realtime;
        filt_in_h_pulse_width 	     			= t_filt_in_h_current_transition - t_filt_in_h_prev_transition;
    end
    else
    begin
        t_filt_in_h_prev_transition 			= 0;
        t_filt_in_h_current_transition 			= 0;
        filt_in_h_pulse_width 				= 0;
    end
end
reg dis_err_msgs;
integer msg_count_pad, msg_count_filt_in_h;
event event_errflag_pad_pulse_width, event_errflag_filt_in_h_pulse_width;
initial
begin
    dis_err_msgs = 1'b1;
    msg_count_pad = 0; msg_count_filt_in_h = 0;


    #1;
    dis_err_msgs = 1'b0;

end
always @(pad_pulse_width)
begin
    if (!dis_err_msgs)
    begin
        if (INP_SEL_H===0 && (pad_pulse_width > min_delay) && (pad_pulse_width < max_delay))
        begin
            msg_count_pad = msg_count_pad + 1;
            ->event_errflag_pad_pulse_width;
            if (msg_count_pad <= MAX_WARNING_COUNT)
            begin
                $display(" ===WARNING=== sky130_fd_io__top_xres4v2 :  Width of Input pulse for PAD input (= %3.2f ns)  is found to be in \the range: %3d ns - %3d ns. In this range, the delay and pulse suppression of the input pulse are PVT dependent. : \%m",pad_pulse_width,min_delay,max_delay,$stime);
            end
            else
                if (msg_count_pad == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_xres4v2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
always @(filt_in_h_pulse_width)
begin
    if (!dis_err_msgs)
    begin
        if (INP_SEL_H===1 && (filt_in_h_pulse_width > min_delay) && (filt_in_h_pulse_width < max_delay))
        begin
            msg_count_filt_in_h = msg_count_filt_in_h + 1;
            ->event_errflag_filt_in_h_pulse_width;
            if (msg_count_filt_in_h <= MAX_WARNING_COUNT)
            begin
                $display(" ===WARNING=== sky130_fd_io__top_xres4v2 :  Width of Input pulse for FILT_IN_H input (= %3.2f ns)  is found to be in \the range: %3d ns - %3d ns. In this range, the delay and pulse suppression of the input pulse are PVT dependent. : \%m",filt_in_h_pulse_width,min_delay,max_delay,$stime);
            end
            else
                if (msg_count_filt_in_h == MAX_WARNING_COUNT+1)
                begin
                    $display(" ===WARNING=== sky130_fd_io__top_xres4v2 :  Further WARNING messages will be suppressed as the \message count has exceeded 100 %m",$stime);
                end
        end
    end
end
endmodule













































































































































































































 // FUNCTIONAL



























































































































































































































































































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_IO__TOP_XRES4V2_V


//--------EOF---------

//-----------------------------------------------------------------------
// Verilog entries for standard power pads (sky130 power pads + overlays)
// Also includes stub entries for the corner and fill cells
// Also includes the custom gpiov2 cell (adds m5 on buses), which is a wrapper
// for the sky130 gpiov2 cell.
//
// This file is distributed as open source under the Apache 2.0 license
// Copyright 2020 efabless, Inc.
// Written by Tim Edwards 
//-----------------------------------------------------------------------

module sky130_ef_io__vccd_hvc_pad (AMUXBUS_A, AMUXBUS_B, DRN_HVC,
	SRC_BDY_HVC, VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VCCD_PAD, VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_HVC;
  inout SRC_BDY_HVC;
  inout VDDIO;	
  inout VDDIO_Q;
  inout VDDA;
  inout VCCD;
  inout VCCD_PAD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD to VCCD)
  sky130_fd_io__top_power_hvc_wpadv2 sky130_fd_io__top_power_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VCCD),
	.P_PAD(VCCD_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(DRN_HVC),
	.SRC_BDY_HVC(SRC_BDY_HVC)
  );

endmodule

module sky130_ef_io__vccd_lvc_pad (AMUXBUS_A, AMUXBUS_B,
	DRN_LVC1, DRN_LVC2, SRC_BDY_LVC1, SRC_BDY_LVC2, BDY2_B2B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VCCD_PAD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_LVC1;
  inout DRN_LVC2;
  inout SRC_BDY_LVC1;
  inout SRC_BDY_LVC2;
  inout BDY2_B2B;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VCCD_PAD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD to VCCD)
  sky130_fd_io__top_power_lvc_wpad sky130_fd_io__top_power_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VCCD),
	.P_PAD(VCCD_PAD),
	.OGC_LVC(),
	.BDY2_B2B(BDY2_B2B),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(DRN_LVC1),
	.DRN_LVC2(DRN_LVC2),
	.SRC_BDY_LVC1(SRC_BDY_LVC1),
	.SRC_BDY_LVC2(SRC_BDY_LVC2)
  );

endmodule

module sky130_ef_io__vdda_lvc_pad (AMUXBUS_A, AMUXBUS_B,
	DRN_LVC1, DRN_LVC2, SRC_BDY_LVC1, SRC_BDY_LVC2, BDY2_B2B,
	VSSA, VDDA, VDDA_PAD, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_LVC1;
  inout DRN_LVC2;
  inout SRC_BDY_LVC1;
  inout SRC_BDY_LVC2;
  inout BDY2_B2B;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VDDA_PAD;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD to VDDA)
  sky130_fd_io__top_power_lvc_wpad sky130_fd_io__top_power_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VDDA),
	.P_PAD(VDDA_PAD),
	.OGC_LVC(),
	.BDY2_B2B(BDY2_B2B),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(DRN_LVC1),
	.DRN_LVC2(DRN_LVC2),
	.SRC_BDY_LVC1(SRC_BDY_LVC1),
	.SRC_BDY_LVC2(SRC_BDY_LVC2)
  );

endmodule

module sky130_ef_io__vdda_hvc_pad (AMUXBUS_A, AMUXBUS_B, DRN_HVC,
	SRC_BDY_HVC,VSSA, VDDA, VDDA_PAD, VSWITCH, VDDIO_Q, VCCHIB,
	VDDIO, VCCD, VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_HVC;
  inout SRC_BDY_HVC;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VDDA_PAD;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD to VDDA)
  sky130_fd_io__top_power_hvc_wpadv2 sky130_fd_io__top_power_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VDDA),
	.P_PAD(VDDA_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(DRN_HVC),
	.SRC_BDY_HVC(SRC_BDY_HVC)
  );

endmodule

module sky130_ef_io__vddio_lvc_pad (AMUXBUS_A, AMUXBUS_B,
	DRN_LVC1, DRN_LVC2, SRC_BDY_LVC1, SRC_BDY_LVC2, BDY2_B2B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VDDIO_PAD, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_LVC1;
  inout DRN_LVC2;
  inout SRC_BDY_LVC1;
  inout SRC_BDY_LVC2;
  inout BDY2_B2B;
  inout VDDIO;	
  inout VDDIO_PAD;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
  sky130_fd_io__top_power_lvc_wpad sky130_fd_io__top_power_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VDDIO),
	.P_PAD(VDDIO_PAD),
	.OGC_LVC(),
	.BDY2_B2B(BDY2_B2B),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(DRN_LVC1),
	.DRN_LVC2(DRN_LVC2),
	.SRC_BDY_LVC1(SRC_BDY_LVC1),
	.SRC_BDY_LVC2(SRC_BDY_LVC2)
  );

  assign VDDIO_Q = VDDIO;

endmodule

module sky130_ef_io__vddio_hvc_pad (AMUXBUS_A, AMUXBUS_B, DRN_HVC,
	SRC_BDY_HVC,VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO,
	VDDIO_PAD, VCCD, VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_HVC;
  inout SRC_BDY_HVC;
  inout VDDIO;	
  inout VDDIO_PAD;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
  sky130_fd_io__top_power_hvc_wpadv2 sky130_fd_io__top_power_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VDDIO),
	.P_PAD(VDDIO_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(DRN_HVC),
	.SRC_BDY_HVC(SRC_BDY_HVC)
  );

  assign VDDIO_Q = VDDIO;

endmodule

module sky130_ef_io__vssd_lvc_pad (AMUXBUS_A, AMUXBUS_B,
	DRN_LVC1, DRN_LVC2, SRC_BDY_LVC1, SRC_BDY_LVC2, BDY2_B2B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSD_PAD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_LVC1;
  inout DRN_LVC2;
  inout SRC_BDY_LVC1;
  inout SRC_BDY_LVC2;
  inout BDY2_B2B;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSD_PAD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying ground pad (connects G_PAD to VSSD)
  sky130_fd_io__top_ground_lvc_wpad sky130_fd_io__top_ground_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSD),
	.G_PAD(VSSD_PAD),
	.OGC_LVC(),
	.BDY2_B2B(BDY2_B2B),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(DRN_LVC1),
	.DRN_LVC2(DRN_LVC2),
	.SRC_BDY_LVC1(SRC_BDY_LVC1),
	.SRC_BDY_LVC2(SRC_BDY_LVC2)
  );

endmodule

module sky130_ef_io__vssd_hvc_pad (AMUXBUS_A, AMUXBUS_B, DRN_HVC,
	SRC_BDY_HVC, VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSD_PAD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_HVC;
  inout SRC_BDY_HVC;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSD_PAD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying ground pad (connects G_PAD to VSSD)
  sky130_fd_io__top_ground_hvc_wpad sky130_fd_io__top_ground_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSD),
	.G_PAD(VSSD_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(DRN_HVC),
	.SRC_BDY_HVC(SRC_BDY_HVC)
  );

endmodule

module sky130_ef_io__vssio_lvc_pad (AMUXBUS_A, AMUXBUS_B,
	DRN_LVC1, DRN_LVC2, SRC_BDY_LVC1, SRC_BDY_LVC2, BDY2_B2B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSIO_PAD, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_LVC1;
  inout DRN_LVC2;
  inout SRC_BDY_LVC1;
  inout SRC_BDY_LVC2;
  inout BDY2_B2B;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;
  inout VSSIO_PAD;

  // Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
  sky130_fd_io__top_ground_lvc_wpad sky130_fd_io__top_ground_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSIO),
	.G_PAD(VSSIO_PAD),
	.OGC_LVC(),
	.BDY2_B2B(BDY2_B2B),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(DRN_LVC1),
	.DRN_LVC2(DRN_LVC2),
	.SRC_BDY_LVC1(SRC_BDY_LVC1),
	.SRC_BDY_LVC2(SRC_BDY_LVC2)
  );

  assign VSSIO_Q = VSSIO;

endmodule


module sky130_ef_io__vssio_hvc_pad (AMUXBUS_A, AMUXBUS_B, DRN_HVC,
	SRC_BDY_HVC,VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSIO_PAD, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_HVC;
  inout SRC_BDY_HVC;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;
  inout VSSIO_PAD;

  // Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
  sky130_fd_io__top_ground_hvc_wpad sky130_fd_io__top_ground_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSIO),
	.G_PAD(VSSIO_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(DRN_HVC),
	.SRC_BDY_HVC(SRC_BDY_HVC)
  );

  assign VSSIO_Q = VSSIO;

endmodule

module sky130_ef_io__vssa_lvc_pad (AMUXBUS_A, AMUXBUS_B,
	DRN_LVC1, DRN_LVC2, SRC_BDY_LVC1, SRC_BDY_LVC2, BDY2_B2B,
	VSSA, VSSA_PAD, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_LVC1;
  inout DRN_LVC2;
  inout SRC_BDY_LVC1;
  inout SRC_BDY_LVC2;
  inout BDY2_B2B;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSA_PAD;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying ground pad (connects G_PAD to VSSA)
  sky130_fd_io__top_ground_lvc_wpad sky130_fd_io__top_ground_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSA),
	.G_PAD(VSSA_PAD),
	.OGC_LVC(),
	.BDY2_B2B(BDY2_B2B),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(DRN_LVC1),
	.DRN_LVC2(DRN_LVC2),
	.SRC_BDY_LVC1(SRC_BDY_LVC1),
	.SRC_BDY_LVC2(SRC_BDY_LVC2)
  );

endmodule

module sky130_ef_io__vssa_hvc_pad (AMUXBUS_A, AMUXBUS_B, DRN_HVC,
	SRC_BDY_HVC,VSSA, VSSA_PAD, VDDA, VSWITCH, VDDIO_Q, VCCHIB,
	VDDIO, VCCD, VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_HVC;
  inout SRC_BDY_HVC;
  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSA_PAD;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying ground pad (connects G_PAD to VSSA)
  sky130_fd_io__top_ground_hvc_wpad sky130_fd_io__top_ground_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSA),
	.G_PAD(VSSA_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(DRN_HVC),
	.SRC_BDY_HVC(SRC_BDY_HVC)
  );

endmodule

module sky130_ef_io__corner_pad (AMUXBUS_A, AMUXBUS_B, 
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

endmodule

module sky130_fd_io__com_bus_slice (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

endmodule

module sky130_ef_io__com_bus_slice_1um (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

endmodule

module sky130_ef_io__com_bus_slice_5um (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

endmodule

module sky130_ef_io__com_bus_slice_10um (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

endmodule

module sky130_ef_io__com_bus_slice_20um (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

endmodule

module sky130_ef_io__gpiov2_pad (IN_H, PAD_A_NOESD_H, PAD_A_ESD_0_H, PAD_A_ESD_1_H,
    PAD, DM, HLD_H_N, IN, INP_DIS, IB_MODE_SEL, ENABLE_H, ENABLE_VDDA_H,
    ENABLE_INP_H, OE_N, TIE_HI_ESD, TIE_LO_ESD, SLOW, VTRIP_SEL, HLD_OVR,
    ANALOG_EN, ANALOG_SEL, ENABLE_VDDIO, ENABLE_VSWITCH_H, ANALOG_POL, OUT,
    AMUXBUS_A, AMUXBUS_B, VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
    VSSIO, VSSD, VSSIO_Q 
    );

input OUT;  		
input OE_N;  		
input HLD_H_N;		
input ENABLE_H;
input ENABLE_INP_H;	
input ENABLE_VDDA_H;	
input ENABLE_VSWITCH_H;	
input ENABLE_VDDIO;	
input INP_DIS;		
input IB_MODE_SEL;
input VTRIP_SEL;	
input SLOW;		
input HLD_OVR;		
input ANALOG_EN;	
input ANALOG_SEL;	
input ANALOG_POL;	
input [2:0] DM;		

inout VDDIO;	
inout VDDIO_Q;	
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;

inout PAD;
inout PAD_A_NOESD_H,PAD_A_ESD_0_H,PAD_A_ESD_1_H;
inout AMUXBUS_A;
inout AMUXBUS_B;

output IN;
output IN_H;
output TIE_HI_ESD, TIE_LO_ESD;

// Instantiate original version with metal4-only power bus
sky130_fd_io__top_gpiov2 gpiov2_base (
    .IN_H(IN_H),
    .PAD_A_NOESD_H(PAD_A_NOESD_H),
    .PAD_A_ESD_0_H(PAD_A_ESD_0_H),
    .PAD_A_ESD_1_H(PAD_A_ESD_1_H),
    .PAD(PAD),
    .DM(DM),
    .HLD_H_N(HLD_H_N),
    .IN(IN),
    .INP_DIS(INP_DIS),
    .IB_MODE_SEL(IB_MODE_SEL),
    .ENABLE_H(ENABLE_H),
    .ENABLE_VDDA_H(ENABLE_VDDA_H),
    .ENABLE_INP_H(ENABLE_INP_H),
    .OE_N(OE_N),
    .TIE_HI_ESD(TIE_HI_ESD),
    .TIE_LO_ESD(TIE_LO_ESD),
    .SLOW(SLOW),
    .VTRIP_SEL(VTRIP_SEL),
    .HLD_OVR(HLD_OVR),
    .ANALOG_EN(ANALOG_EN),
    .ANALOG_SEL(ANALOG_SEL),
    .ENABLE_VDDIO(ENABLE_VDDIO),
    .ENABLE_VSWITCH_H(ENABLE_VSWITCH_H),
    .ANALOG_POL(ANALOG_POL),
    .OUT(OUT),
    .AMUXBUS_A(AMUXBUS_A),
    .AMUXBUS_B(AMUXBUS_B),
    .VSSA(VSSA),
    .VDDA(VDDA),
    .VSWITCH(VSWITCH),
    .VDDIO_Q(VDDIO_Q),
    .VCCHIB(VCCHIB),
    .VDDIO(VDDIO),
    .VCCD(VCCD),
    .VSSIO(VSSIO),
    .VSSD(VSSD),
    .VSSIO_Q(VSSIO_Q) 
);

endmodule

// sky130_ef_io__vddio_hvc_pad with HV clamp connections to VDDIO and VSSIO

module sky130_ef_io__vddio_hvc_clamped_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VDDIO_PAD, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;
  inout VDDIO_PAD;
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
  sky130_fd_io__top_power_hvc_wpadv2 sky130_fd_io__top_power_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VDDIO),
	.P_PAD(VDDIO_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(VDDIO),
	.SRC_BDY_HVC(VSSIO)
  );

  assign VDDIO_Q = VDDIO;

endmodule

// sky130_ef_io__vssio_hvc_pad with HV clamp connections to VDDIO and VSSIO

module sky130_ef_io__vssio_hvc_clamped_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSIO_PAD, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;
  inout VSSIO_PAD;

  // Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
  sky130_fd_io__top_ground_hvc_wpad sky130_fd_io__top_ground_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSIO),
	.G_PAD(VSSIO_PAD),
	.OGC_HVC(VDDIO),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(VDDIO),
	.SRC_BDY_HVC(VSSIO)
  );

  assign VSSIO_Q = VSSIO;

endmodule

// sky130_ef_io__vdda_hvc_pad with HV clamp connections to VDDA and VSSA

module sky130_ef_io__vdda_hvc_clamped_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VDDA_PAD, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VDDA_PAD;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD to VDDA)
  sky130_fd_io__top_power_hvc_wpadv2 sky130_fd_io__top_power_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VDDA),
	.P_PAD(VDDA_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(VDDA),
	.SRC_BDY_HVC(VSSA)
  );

endmodule

// sky130_ef_io__vssa_hvc_pad with HV clamp connections to VDDA and VSSA

module sky130_ef_io__vssa_hvc_clamped_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VSSA_PAD, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSA_PAD;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying ground pad (connects G_PAD to VSSA)
  sky130_fd_io__top_ground_hvc_wpad sky130_fd_io__top_ground_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSA),
	.G_PAD(VSSA_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(VDDA),
	.SRC_BDY_HVC(VSSA)
  );

endmodule

// sky130_ef_io__vccd_lvc_pad with LV clamp connections to VCCD/VSSIO and VCCD/VSSD,
// and back-to-back diodes connecting VSSIO to VSSA

module sky130_ef_io__vccd_lvc_clamped_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VCCD_PAD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VCCD_PAD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD to VCCD)
  sky130_fd_io__top_power_lvc_wpad sky130_fd_io__top_power_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VCCD),
	.P_PAD(VCCD_PAD),
	.OGC_LVC(),
	.BDY2_B2B(VSSA),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(VCCD),
	.DRN_LVC2(VCCD),
	.SRC_BDY_LVC1(VSSIO),
	.SRC_BDY_LVC2(VSSD)
  );

endmodule

// sky130_ef_io__vssd_lvc_pad with LV clamp connections to VCCD/VSSIO and VCCD/VSSD,
// and back-to-back diodes connecting VSSIO to VSSA

module sky130_ef_io__vssd_lvc_clamped_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSD_PAD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSD_PAD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying ground pad (connects G_PAD to VSSD)
  sky130_fd_io__top_ground_lvc_wpad sky130_fd_io__top_ground_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSD),
	.G_PAD(VSSD_PAD),
	.OGC_LVC(),
	.BDY2_B2B(VSSA),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(VCCD),
	.DRN_LVC2(VCCD),
	.SRC_BDY_LVC1(VSSIO),
	.SRC_BDY_LVC2(VSSD)
  );

endmodule

// sky130_ef_io__vccd_lvc_pad with LV clamp connections to VCCD and VSSD,
// and back-to-back diodes connecting VSSD to VSSIO

module sky130_ef_io__vccd_lvc_clamped2_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VCCD_PAD,
	VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VCCD_PAD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD to VCCD)
  sky130_fd_io__top_power_lvc_wpad sky130_fd_io__top_power_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VCCD),
	.P_PAD(VCCD_PAD),
	.OGC_LVC(),
	.BDY2_B2B(VSSIO),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(VCCD),
	.DRN_LVC2(VCCD),
	.SRC_BDY_LVC1(VSSD),
	.SRC_BDY_LVC2(VSSD)
  );

endmodule

// sky130_ef_io__vssd_lvc_pad with LV clamp connections to VCCD and VSSD,
// and back-to-back diodes connecting VSSD to VSSIO

module sky130_ef_io__vssd_lvc_clamped2_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSD_PAD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSD_PAD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying ground pad (connects G_PAD to VSSD)
  sky130_fd_io__top_ground_lvc_wpad sky130_fd_io__top_ground_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSD),
	.G_PAD(VSSD_PAD),
	.OGC_LVC(),
	.BDY2_B2B(VSSIO),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(VCCD),
	.DRN_LVC2(VCCD),
	.SRC_BDY_LVC1(VSSD),
	.SRC_BDY_LVC2(VSSD)
  );

endmodule

// sky130_ef_io__vccd_lvc_pad with pad and LV clamp connection to VCCD1,
// pad negative connection to VSSD1, and back-to-back diodes connecting
// VSSD1 to VSSIO

module sky130_ef_io__vccd_lvc_clamped3_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD, VCCD_PAD,
	VSSIO, VSSD, VSSIO_Q, VCCD1, VSSD1
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VCCD_PAD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;
  inout VCCD1;
  inout VSSD1;

  // Instantiate the underlying power pad (connects P_PAD to VCCD1)
  sky130_fd_io__top_power_lvc_wpad sky130_fd_io__top_power_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(VCCD1),
	.P_PAD(VCCD_PAD),
	.OGC_LVC(),
	.BDY2_B2B(VSSIO),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(VCCD1),
	.DRN_LVC2(VCCD1),
	.SRC_BDY_LVC1(VSSD1),
	.SRC_BDY_LVC2(VSSD1)
  );

endmodule

// sky130_ef_io__vssd_lvc_pad with pad and LV clamp negative connection
// to VSSD1, clamp positive connection to VCCD1, and back-to-back diodes
// connecting VSSD1 to VSSIO

module sky130_ef_io__vssd_lvc_clamped3_pad (AMUXBUS_A, AMUXBUS_B,
	VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
	VSSIO, VSSD, VSSD_PAD, VSSIO_Q, VCCD1, VSSD1
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout VDDIO;	
  inout VDDIO_Q;	
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSD_PAD;
  inout VSSIO_Q;
  inout VSSIO;
  inout VCCD1;
  inout VSSD1;

  // Instantiate the underlying ground pad (connects G_PAD to VSSD1)
  sky130_fd_io__top_ground_lvc_wpad sky130_fd_io__top_ground_lvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.G_CORE(VSSD1),
	.G_PAD(VSSD_PAD),
	.OGC_LVC(),
	.BDY2_B2B(VSSIO),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_LVC1(VCCD1),
	.DRN_LVC2(VCCD1),
	.SRC_BDY_LVC1(VSSD1),
	.SRC_BDY_LVC2(VSSD1)
  );

endmodule

// 

module sky130_ef_io__top_power_hvc (AMUXBUS_A, AMUXBUS_B, DRN_HVC,
	P_CORE, P_PAD, SRC_BDY_HVC, VSSA, VDDA, VSWITCH, VDDIO_Q,
	VCCHIB, VDDIO, VCCD, VSSIO, VSSD, VSSIO_Q
);
  inout AMUXBUS_A;
  inout AMUXBUS_B;

  inout DRN_HVC;
  inout P_CORE;
  inout P_PAD;
  inout SRC_BDY_HVC;
  inout VDDIO;	
  inout VDDIO_Q;
  inout VDDA;
  inout VCCD;
  inout VSWITCH;
  inout VCCHIB;
  inout VSSA;
  inout VSSD;
  inout VSSIO_Q;
  inout VSSIO;

  // Instantiate the underlying power pad (connects P_PAD to VCCD)
  sky130_fd_io__top_power_hvc_wpadv2 sky130_fd_io__top_power_hvc_base ( 
	.VSSA(VSSA),
	.VDDA(VDDA),
	.VSWITCH(VSWITCH),
	.VDDIO_Q(VDDIO_Q),
	.VCCHIB(VCCHIB),
	.VDDIO(VDDIO),
	.VCCD(VCCD),
	.VSSIO(VSSIO),
	.VSSD(VSSD),
	.VSSIO_Q(VSSIO_Q),
	.P_CORE(P_CORE),
	.P_PAD(P_PAD),
	.OGC_HVC(),
	.AMUXBUS_A(AMUXBUS_A),
	.AMUXBUS_B(AMUXBUS_B),
	.DRN_HVC(DRN_HVC),
	.SRC_BDY_HVC(SRC_BDY_HVC)
  );

endmodule



//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * analog_pad: Analog PAD.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none





/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/

module sky130_ef_io__analog_pad (AMUXBUS_A, AMUXBUS_B, P_PAD, P_CORE
                                 ,VCCD, VCCHIB, VDDA, VDDIO, VDDIO_Q, VSSA, VSSD, VSSIO, VSSIO_Q, VSWITCH
                                );
inout AMUXBUS_A;
inout AMUXBUS_B;
inout P_PAD;
inout P_CORE;
inout VCCD;
inout VCCHIB;
inout VDDA;
inout VDDIO;
inout VDDIO_Q;
inout VSSA;
inout VSSD;
inout VSSIO;
inout VSSIO_Q;
inout VSWITCH;
wire pwr_good = VDDIO===1 && VSSIO===0;
wire pad_sw = pwr_good===1 ? 1'b1 : 1'bx;
tranif1 x_pad (P_PAD, P_CORE, pad_sw);
endmodule











































 // FUNCTIONAL























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_EF_IO__ANALOG_PAD_V


//--------EOF---------

module sky130_ef_io__gpiov2_pad_wrapped (IN_H, PAD_A_NOESD_H, PAD_A_ESD_0_H, PAD_A_ESD_1_H,
    PAD, DM, HLD_H_N, IN, INP_DIS, IB_MODE_SEL, ENABLE_H, ENABLE_VDDA_H,
    ENABLE_INP_H, OE_N, TIE_HI_ESD, TIE_LO_ESD, SLOW, VTRIP_SEL, HLD_OVR,
    ANALOG_EN, ANALOG_SEL, ENABLE_VDDIO, ENABLE_VSWITCH_H, ANALOG_POL, OUT,
    AMUXBUS_A, AMUXBUS_B, VSSA, VDDA, VSWITCH, VDDIO_Q, VCCHIB, VDDIO, VCCD,
    VSSIO, VSSD, VSSIO_Q 
    );

input OUT;  		
input OE_N;  		
input HLD_H_N;		
input ENABLE_H;
input ENABLE_INP_H;	
input ENABLE_VDDA_H;	
input ENABLE_VSWITCH_H;	
input ENABLE_VDDIO;	
input INP_DIS;		
input IB_MODE_SEL;
input VTRIP_SEL;	
input SLOW;		
input HLD_OVR;		
input ANALOG_EN;	
input ANALOG_SEL;	
input ANALOG_POL;	
input [2:0] DM;		

inout VDDIO;	
inout VDDIO_Q;	
inout VDDA;
inout VCCD;
inout VSWITCH;
inout VCCHIB;
inout VSSA;
inout VSSD;
inout VSSIO_Q;
inout VSSIO;

inout PAD;
inout PAD_A_NOESD_H,PAD_A_ESD_0_H,PAD_A_ESD_1_H;
inout AMUXBUS_A;
inout AMUXBUS_B;

output IN;
output IN_H;
output TIE_HI_ESD, TIE_LO_ESD;

// Instantiate original version with metal4-only power bus
sky130_fd_io__top_gpiov2 gpiov2_base (
    .IN_H(IN_H),
    .PAD_A_NOESD_H(PAD_A_NOESD_H),
    .PAD_A_ESD_0_H(PAD_A_ESD_0_H),
    .PAD_A_ESD_1_H(PAD_A_ESD_1_H),
    .PAD(PAD),
    .DM(DM),
    .HLD_H_N(HLD_H_N),
    .IN(IN),
    .INP_DIS(INP_DIS),
    .IB_MODE_SEL(IB_MODE_SEL),
    .ENABLE_H(ENABLE_H),
    .ENABLE_VDDA_H(ENABLE_VDDA_H),
    .ENABLE_INP_H(ENABLE_INP_H),
    .OE_N(OE_N),
    .TIE_HI_ESD(TIE_HI_ESD),
    .TIE_LO_ESD(TIE_LO_ESD),
    .SLOW(SLOW),
    .VTRIP_SEL(VTRIP_SEL),
    .HLD_OVR(HLD_OVR),
    .ANALOG_EN(ANALOG_EN),
    .ANALOG_SEL(ANALOG_SEL),
    .ENABLE_VDDIO(ENABLE_VDDIO),
    .ENABLE_VSWITCH_H(ENABLE_VSWITCH_H),
    .ANALOG_POL(ANALOG_POL),
    .OUT(OUT),
    .AMUXBUS_A(AMUXBUS_A),
    .AMUXBUS_B(AMUXBUS_B),
    .VSSA(VSSA),
    .VDDA(VDDA),
    .VSWITCH(VSWITCH),
    .VDDIO_Q(VDDIO_Q),
    .VCCHIB(VCCHIB),
    .VDDIO(VDDIO),
    .VCCD(VCCD),
    .VSSIO(VSSIO),
    .VSSD(VSSD),
    .VSSIO_Q(VSSIO_Q) 
);

endmodule


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog wrapper for decap with size of 12 units.
 * This cell has been modified from sky130_fd_sc_hd__decap_12
 * to remove excess LI, so that when used extensively in a
 * padded region of a digital layout, it does not cause the
 * LI layer to exceed critical density.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_ef_sc_hd__decap_12 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__decap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_EF_SC_HD__DECAP_12_V




//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fakediode: Antenna tie-down diode with no connection between the DIODE
 * pin and the diode.  This is just the sky130_fd_sc_hd__diode_2 cell with
 * the contacts removed between the diode and the pin.  It is used by the
 * openlane synthesis flow to preemptively put antenna tie-downs close to
 * every pin without making a connection.  If the net needs an antenna
 * tiedown, the fakediode cell can be replaced by the real diode cell.
 *
 * Verilog wrapper for diode with size of 2 units.  Note that the wrapper
 * is around the original SkyWater diode base cell;  because the diode
 * has no function in verilog, there is no difference between the verilog
 * definitions of the diode and fake diode other than the cell name.
 *
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_ef_sc_hd__fakediode_2 (
    DIODE,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    input DIODE;
    input VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__diode base (
        .DIODE(DIODE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/
























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_EF_SC_HD__FAKEDIODE_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none


/*********************************************************/

`celldefine
module sky130_ef_sc_hd__fill_8 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;

endmodule
`endcelldefine

/*********************************************************/















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_EF_SC_HD__FILL_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill_12:  Designed to replace the decap_12 cell while reducing the
 * amount of local interconnect;  this is just a decap_6, fill_4, and
 * fill_2 cell juxtaposed, making up the same width as the decap_12
 * but with half the amount of decap.
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_ef_sc_hd__fill_12 (
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    input VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_EF_SC_HD__FILL_12_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$NSR: Negative edge triggered D flip-flop (Q output UDP)
 *              with both active high reset and set (set dominate).
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dff$NSR (
    Q    ,
    SET  ,
    RESET,
    CLK_N,
    D
);

    output Q    ;
    input  SET  ;
    input  RESET;
    input  CLK_N;
    input  D    ;

    reg Q;

    table
     // SET RESET CLK_N  D  :  Qt : Qt+1
         0    1     ?    ?  :  ?  :  0    ; // Asserting reset
         0    *     ?    ?  :  0  :  0    ; // Changing reset
         1    ?     ?    ?  :  ?  :  1    ; // Asserting set (dominates reset)
         *    0     ?    ?  :  1  :  1    ; // Changing set
         0    ?    (01)  0  :  ?  :  0    ; // rising clock
         ?    0    (01)  1  :  ?  :  1    ; // rising clock
         0    ?     p    0  :  0  :  0    ; // potential rising clock
         ?    0     p    1  :  1  :  1    ; // potential rising clock
         0    0     n    ?  :  ?  :  -    ; // Clock falling register output does not change
         0    0     ?    *  :  ?  :  -    ; // Changing Data
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DFF_NSR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$NSR_pp$PG$N: Negative edge triggered D flip-flop
 *                      (Q output UDP) with both active high reset and
 *                      set (set dominate). Includes VPWR and VGND
 *                      power pins and notifier pin.
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dff$NSR_pp$PG$N (
    Q       ,
    SET     ,
    RESET   ,
    CLK_N   ,
    D       ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  SET     ;
    input  RESET   ;
    input  CLK_N   ;
    input  D       ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //         SET          RESET CLK_N  D  NOTIFIER VPWR VGND :  Qt : Qt+1
                 0             1     b    ?     ?      1    0   :  ?  :  0    ; // Asserting reset
                 0             *     ?    ?     ?      1    0   :  0  :  0    ; // Changing reset
                 1             ?     b    ?     ?      1    0   :  ?  :  1    ; // Asserting set  (dominates reset)
                 *             0     ?    ?     ?      1    0   :  1  :  1    ; // Changing set
                 1             ?     n    ?     ?      1    0   :  1  :  1    ;
                 ?             1     n    ?     ?      1    0   :  0  :  0    ;
                 x             ?     n    ?     ?      1    0   :  1  :  1    ;
                 ?             x     n    ?     ?      1    0   :  0  :  0    ;
                 0             ?    (01)  0     ?      1    0   :  ?  :  0    ; // rising clock
                 ?             0    (01)  1     ?      1    0   :  ?  :  1    ; // rising clock
                 0             ?     p    0     ?      1    0   :  0  :  0    ; // potential rising clock
                 ?             0     p    1     ?      1    0   :  1  :  1    ; // potential rising clock
                 0             ?     x    0     ?      1    0   :  1  :  x    ;
                 ?             0     x    1     ?      1    0   :  0  :  x    ;
                 0             0     n    ?     ?      1    0   :  ?  :  -    ; // Clock falling register output does not change
                 0             0     ?    *     ?      1    0   :  ?  :  -    ; // Changing Data
        // ['IfDef(functional)', '']                 ?             ?     ?    ?     *      1    0   :  ?  :  -    ; // go to - on notify
        // ['Else', '']                 ?             ?     ?    ?     *      1    0   :  ?  :  X    ; // go to X on notify
        // ['EndIfDef(functional)', '']                 ?             ?     ?    ?     ?      *    0   :  ?  :  X    ; // any change on vpwr
                 ?             ?     ?    ?     ?      ?    *   :  ?  :  X    ; // any change on vgnd
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DFF_NSR_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$P: Positive edge triggered D flip-flop (Q output UDP).
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dff$P (
    Q  ,
    D  ,
    CLK
);

    output Q  ;
    input  D  ;
    input  CLK;

    reg Q;

    table
     //  D  CLK  :  Qt : Qt+1
         1  (01) :  ?  :  1    ; // clocked data
         0  (01) :  ?  :  0    ;
         1  (x1) :  1  :  1    ; // reducing pessimism
         0  (x1) :  0  :  0    ;
         1  (0x) :  1  :  1    ;
         0  (0x) :  0  :  0    ;
         ?  (1x) :  ?  :  -    ; // no change on falling edge
         ?  (?0) :  ?  :  -    ;
         *   ?   :  ?  :  -    ; // ignore edges on data
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DFF_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$P_pp$PG$N: Positive edge triggered D flip-flop
 *                    (Q output UDP).
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dff$P_pp$PG$N (
    Q       ,
    D       ,
    CLK     ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  CLK     ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           CLK  NOTIFIER VPWR VGND :  Qt : Qt+1
                 1           (01)    ?      1    0   :  ?  :  1    ; // clocked data
                 0           (01)    ?      1    0   :  ?  :  0    ;
                 1           (x1)    ?      1    0   :  1  :  1    ; // reducing pessimism
                 0           (x1)    ?      1    0   :  0  :  0    ;
                 1           (0x)    ?      1    0   :  1  :  1    ;
                 0           (0x)    ?      1    0   :  0  :  0    ;
                 0            x      ?      1    0   :  0  :  0    ; // Hold when CLK=X and D=Q
                 1            x      ?      1    0   :  1  :  1    ; // Hold when CLK=X and D=Q
                 ?           (?0)    ?      1    0   :  ?  :  -    ;
                 *            b      ?      1    0   :  ?  :  -    ; // ignore edges on data
        // ['IfDef(functional)', '']                 ?            ?      *      1    0   :  ?  :  -    ;
        // ['Else', '']                 ?            ?      *      1    0   :  ?  :  x    ;
        // ['EndIfDef(functional)', '']                 ?            ?      ?      *    ?   :  ?  :  x    ; // any change on vpwr
                 ?            ?      ?      ?    *   :  ?  :  x    ; // any change on vgnd
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DFF_P_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$PR: Positive edge triggered D flip-flop with active high
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dff$PR (
    Q    ,
    D    ,
    CLK  ,
    RESET
);

    output Q    ;
    input  D    ;
    input  CLK  ;
    input  RESET;

    reg Q;

    table
     //  D  CLK  RESET :  Qt : Qt+1
         *   b     0   :  ?  :  -    ; // data event, hold unless CP==x
         ?  (?0)   0   :  ?  :  -    ; // CP => 0, hold
         ?   b    (?0) :  ?  :  -    ; // R => 0, hold unless CP==x
         ?   ?     1   :  ?  :  0    ; // async reset
         0   r     ?   :  ?  :  0    ; // clock data on CP
         1   r     0   :  ?  :  1    ; // clock data on CP
         0  (x1)   ?   :  0  :  0    ; // possible CP, hold when D==Q==0
         1  (x1)   0   :  1  :  1    ; // possible CP, hold when D==Q==1
         0   x     ?   :  0  :  0    ; // unkown CP, hold when D==Q==0
         1   x     0   :  1  :  1    ; // unkown CP, hold when D==Q==1
         ?   b    (?x) :  0  :  0    ; // R=>x, hold when Q==0 unless CP==x
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DFF_PR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$PR_pp$PG$N: Positive edge triggered D flip-flop with active
 *                     high
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dff$PR_pp$PG$N (
    Q       ,
    D       ,
    CLK     ,
    RESET   ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  CLK     ;
    input  RESET   ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           CLK  RESET NOTIFIER VPWR VGND :  Qt : Qt+1
                 *            b     0      ?      1    0   :  ?  :  -    ; // data event, hold unless CP==x
                 ?           (?0)   0      ?      1    0   :  ?  :  -    ; // CP => 0, hold
                 ?            b    (?0)    ?      1    0   :  ?  :  -    ; // R => 0, hold unless CP==x
                 ?            ?     1      ?      1    0   :  ?  :  0    ; // async reset
                 0            r     ?      ?      1    0   :  ?  :  0    ; // clock data on CP
                 1            r     0      ?      1    0   :  ?  :  1    ; // clock data on CP
                 0           (x1)   ?      ?      1    0   :  0  :  0    ; // possible CP, hold when D==Q==0
                 1           (x1)   0      ?      1    0   :  1  :  1    ; // possible CP, hold when D==Q==1
                 0            x     ?      ?      1    0   :  0  :  0    ; // unkown CP, hold when D==Q==0
                 1            x     0      ?      1    0   :  1  :  1    ; // unkown CP, hold when D==Q==1
                 ?            b    (?x)    ?      1    0   :  0  :  0    ; // R=>x, hold when Q==0 unless CP==x
                 ?           (?0)   x      ?      1    0   :  0  :  0    ;
        // ['IfDef(functional)', '']                 ?            ?     ?      *      1    0   :  ?  :  -    ; // Q => - on any change on notifier
        // ['Else', '']                 ?            ?     ?      *      1    0   :  ?  :  x    ; // Q => X on any change on notifier
        // ['EndIfDef(functional)', '']                 ?            ?     ?      ?      *    ?   :  ?  :  x    ; // Q => X on any change on vpwr
                 ?            ?     ?      ?      ?    *   :  ?  :  x    ; // Q => X on any change on vgnd
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DFF_PR_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$PS: Positive edge triggered D flip-flop with active high
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dff$PS (
    Q  ,
    D  ,
    CLK,
    SET
);

    output Q  ;
    input  D  ;
    input  CLK;
    input  SET;

    reg Q;

    table
     //  D  CLK  SET  :  Qt : Qt+1
         *   b    0   :  ?  :  -    ; // data event, hold unless CP==x
         ?  (?0)  0   :  ?  :  -    ; // CP => 0, hold
         ?   b   (?0) :  ?  :  -    ; // S => 0, hold unless CP==x
         ?   ?    1   :  ?  :  1    ; // async set
         0   r    0   :  ?  :  0    ; // clock data on CP
         1   r    ?   :  ?  :  1    ; // clock data on CP
         0  (x1)  0   :  0  :  0    ; // possible CP, hold when D==Q==0
         1  (x1)  ?   :  1  :  1    ; // possible CP, hold when D==Q==1
         0   x    0   :  0  :  0    ; // unkown CP, hold when D==Q==0
         1   x    ?   :  1  :  1    ; // unkown CP, hold when D==Q==1
         ?   b   (?x) :  1  :  1    ; // S=>x, hold when Q==1 unless CP==x
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DFF_PS_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$PS_pp$PG$N: Positive edge triggered D flip-flop with active
 *                     high
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dff$PS_pp$PG$N (
    Q       ,
    D       ,
    CLK     ,
    SET     ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  CLK     ;
    input  SET     ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           CLK  SET  NOTIFIER VPWR VGND :  Qt : Qt+1
                 *            b    0      ?      1    0   :  ?  :  -    ; // data event, hold unless CP==x
                 ?           (?0)  0      ?      1    0   :  ?  :  -    ; // CP => 0, hold
                 ?            b   (?0)    ?      1    0   :  ?  :  -    ; // S => 0, hold unless CP==x
                 ?            ?    1      ?      1    0   :  ?  :  1    ; // async set
                 0            r    0      ?      1    0   :  ?  :  0    ; // clock data on CP
                 1            r    ?      ?      1    0   :  ?  :  1    ; // clock data on CP
                 0           (x1)  0      ?      1    0   :  0  :  0    ; // possible CP, hold when D==Q==0
                 1           (x1)  ?      ?      1    0   :  1  :  1    ; // possible CP, hold when D==Q==1
                 0            x    0      ?      1    0   :  0  :  0    ; // unkown CP, hold when D==Q==0
                 1            x    ?      ?      1    0   :  1  :  1    ; // unkown CP, hold when D==Q==1
                 ?            b   (?x)    ?      1    0   :  1  :  1    ; // S=>x, hold when Q==1 unless CP==x
                 ?           (?0)  x      ?      1    0   :  1  :  1    ;
        // ['IfDef(functional)', '']                 ?            ?    ?      *      1    0   :  ?  :  -    ; // Q => - on any change on notifier
        // ['Else', '']                 ?            ?    ?      *      1    0   :  ?  :  x    ; // Q => X on any change on notifier
        // ['EndIfDef(functional)', '']                 ?            ?    ?      ?      *    ?   :  ?  :  x    ; // Q => X on any change on vpwr
                 ?            ?    ?      ?      ?    *   :  ?  :  x    ; // Q => X on any change on vgnd
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DFF_PS_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$lP: D-latch, gated standard drive / active high
 *                (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dlatch$lP (
    Q   ,
    D   ,
    GATE
);

    output Q   ;
    input  D   ;
    input  GATE;

    reg Q;

    table
     //  D  GATE :  Qt : Qt+1
         ?   0   :  ?  :  -    ; // hold
         0   1   :  ?  :  0    ; // pass 0
         1   1   :  ?  :  1    ; // pass 1
         0   x   :  0  :  0    ; // reduce pessimism
         1   x   :  1  :  1    ; // reduce pessimism
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DLATCH_LP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$lP_pp$PG$N: D-latch, gated standard drive / active high
 *                        (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dlatch$lP_pp$PG$N (
    Q       ,
    D       ,
    GATE    ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  GATE    ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           GATE NOTIFIER VPWR VGND : Qtn : Qtn+1
                 *            0      ?      1    0   :  ?  :   -    ;
                 ?           (?0)    ?      1    0   :  ?  :   -    ;
                 ?           (1x)    ?      1    0   :  ?  :   -    ;
                 0           (0x)    ?      1    0   :  0  :   0    ;
                 1           (0x)    ?      1    0   :  1  :   1    ;
                 0           (x1)    ?      1    0   :  ?  :   0    ;
                 1           (x1)    ?      1    0   :  ?  :   1    ;
                (?0)          1      ?      1    0   :  ?  :   0    ;
                (?1)          1      ?      1    0   :  ?  :   1    ;
                 0           (01)    ?      1    0   :  ?  :   0    ;
                 1           (01)    ?      1    0   :  ?  :   1    ;
                (?1)          x      ?      1    0   :  1  :   1    ; // Reducing pessimism.
                (?0)          x      ?      1    0   :  0  :   0    ;
        // ['IfDef(functional)', '']                 ?            ?      *      1    0   :  ?  :   -    ;
        // ['Else', '']                 ?            ?      *      1    0   :  ?  :   x    ;
        // ['EndIfDef(functional)', '']                 ?            ?      ?      *    ?   :  ?  :   x    ; // any change on vpwr
                 ?            ?      ?      ?    *   :  ?  :   x    ; // any change on vgnd
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DLATCH_LP_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$P: D-latch, gated standard drive / active high
 *               (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dlatch$P (
    Q   ,
    D   ,
    GATE
);

    output Q   ;
    input  D   ;
    input  GATE;

    reg Q;

    table
     //  D  GATE :  Qt : Qt+1
         ?   0   :  ?  :  -    ; // hold
         0   1   :  ?  :  0    ; // pass 0
         1   1   :  ?  :  1    ; // pass 1
         0   x   :  0  :  0    ; // reduce pessimism
         1   x   :  1  :  1    ; // reduce pessimism
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DLATCH_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$P_pp$PG$N: D-latch, gated standard drive / active high
 *                       (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dlatch$P_pp$PG$N (
    Q       ,
    D       ,
    GATE    ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  GATE    ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           GATE NOTIFIER VPWR VGND : Qtn : Qtn+1
                 *            0      ?      1    0   :  ?  :   -    ;
                 ?           (?0)    ?      1    0   :  ?  :   -    ;
                 ?           (1x)    ?      1    0   :  ?  :   -    ;
                 0           (0x)    ?      1    0   :  0  :   0    ;
                 1           (0x)    ?      1    0   :  1  :   1    ;
                 0           (x1)    ?      1    0   :  ?  :   0    ;
                 1           (x1)    ?      1    0   :  ?  :   1    ;
                (?0)          1      ?      1    0   :  ?  :   0    ;
                (?1)          1      ?      1    0   :  ?  :   1    ;
                 0           (01)    ?      1    0   :  ?  :   0    ;
                 1           (01)    ?      1    0   :  ?  :   1    ;
                (?1)          x      ?      1    0   :  1  :   1    ; // Reducing pessimism.
                (?0)          x      ?      1    0   :  0  :   0    ;
        // ['IfDef(functional)', '']                 ?            ?      *      1    0   :  ?  :   -    ;
        // ['Else', '']                 ?            ?      *      1    0   :  ?  :   x    ;
        // ['EndIfDef(functional)', '']                 0            1      ?     (?1)  0   :  ?  :   0    ;
                 1            1      ?     (?1)  0   :  ?  :   1    ;
                 0            1      ?      1   (?0) :  ?  :   0    ;
                 1            1      ?      1   (?0) :  ?  :   1    ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DLATCH_P_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$PR: D-latch, gated clear direct / gate active high
 *                (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dlatch$PR (
    Q    ,
    D    ,
    GATE ,
    RESET
);

    output Q    ;
    input  D    ;
    input  GATE ;
    input  RESET;

    reg Q;

    table
     //  D  GATE RESET :  Qt : Qt+1
         ?   0     0   :  ?  :  -    ; // hold
         0   1     0   :  ?  :  0    ; // pass 0
         1   1     0   :  ?  :  1    ; // pass 1
         ?   ?     1   :  ?  :  0    ; // async reset
         0   1     ?   :  ?  :  0    ; // reduce pessimism
         0   x     0   :  0  :  0    ; // reduce pessimism
         1   x     0   :  1  :  1    ; // reduce pessimism
         ?   0     x   :  0  :  0    ; // reduce pessimism
         0   x     x   :  0  :  0    ; // reduce pessimism
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DLATCH_PR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$PR_pp$PG$N: D-latch, gated clear direct / gate active
 *                        high (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_dlatch$PR_pp$PG$N (
    Q       ,
    D       ,
    GATE    ,
    RESET   ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  GATE    ;
    input  RESET   ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           GATE RESET NOTIFIER VPWR VGND :  Qt : Qt+1
                 *            0     0      ?      1    0   :  ?  :  -    ;
                 ?            ?     1      ?      1    0   :  ?  :  0    ; // asynchro clear
                 ?           (?0)   0      ?      1    0   :  ?  :  -    ; // Changed R=? to R=0 ; jek 08/14/06/
                 ?           (1x)   0      ?      1    0   :  ?  :  -    ; // Changed R=? to R=0 ; jek 08/14/06
                 0           (0x)   0      ?      1    0   :  0  :  0    ;
                 1           (0x)   0      ?      1    0   :  1  :  1    ;
                 0           (x1)   0      ?      1    0   :  ?  :  0    ;
                 1           (x1)   0      ?      1    0   :  ?  :  1    ;
                (?0)          1     0      ?      1    0   :  ?  :  0    ;
                (?1)          1     0      ?      1    0   :  ?  :  1    ;
                 0           (01)   0      ?      1    0   :  ?  :  0    ;
                 1           (01)   0      ?      1    0   :  ?  :  1    ;
                 ?            0    (?x)    ?      1    0   :  0  :  0    ; // Reducing pessimism.//AB
                 *            0     x      ?      1    0   :  0  :  0    ; // Reducing pessimism//AB
                 0           (?1)   x      ?      1    0   :  ?  :  0    ; // Reducing pessimism.
                (?0)          1     x      ?      1    0   :  ?  :  0    ; // Reducing pessimism.
                 0            1    (?x)    ?      1    0   :  ?  :  0    ; // Reducing pessimism.//AB
                 ?            0    (?0)    ?      1    0   :  ?  :  -    ; // ignore edge on clear
                 0            1    (?0)    ?      1    0   :  ?  :  0    ; // pessimism .
                 1            1    (?0)    ?      1    0   :  ?  :  1    ;
                (?1)          x     0      ?      1    0   :  1  :  1    ; // Reducing pessimism.
                (?0)          x     0      ?      1    0   :  0  :  0    ; // Reducing pessimism.
        // ['IfDef(functional)', '']                 ?            ?     ?      *      1    0   :  ?  :  -    ;
        // ['Else', '']                 ?            ?     ?      *      1    0   :  ?  :  x    ;
        // ['EndIfDef(functional)', '']                 0            1     0      ?     (?1)  0   :  ?  :  0    ;
                 1            1     0      ?     (?1)  0   :  ?  :  1    ;
                 0            1     0      ?      1   (?0) :  ?  :  0    ;
                 1            1     0      ?      1   (?0) :  ?  :  1    ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_DLATCH_PR_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_mux_2to1: Two to one multiplexer
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_mux_2to1 (
    X ,
    A0,
    A1,
    S
);

    output X ;
    input  A0;
    input  A1;
    input  S ;

    table
     //  A0  A1  S  :  X
         0   0   ?  :  0   ;
         1   1   ?  :  1   ;
         0   ?   0  :  0   ;
         1   ?   0  :  1   ;
         ?   0   1  :  0   ;
         ?   1   1  :  1   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_MUX_2TO1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_mux_2to1_N: Two to one multiplexer with inverting output
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_mux_2to1_N (
    Y ,
    A0,
    A1,
    S
);

    output Y ;
    input  A0;
    input  A1;
    input  S ;

    table
     //  A0  A1  S  :  Y
         0   ?   0  :  1   ;
         1   ?   0  :  0   ;
         ?   0   1  :  1   ;
         ?   1   1  :  0   ;
         0   0   ?  :  1   ;
         1   1   ?  :  0   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_MUX_2TO1_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_mux_4to2: Four to one multiplexer with 2 select controls
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_mux_4to2 (
    X ,
    A0,
    A1,
    A2,
    A3,
    S0,
    S1
);

    output X ;
    input  A0;
    input  A1;
    input  A2;
    input  A3;
    input  S0;
    input  S1;

    table
     //  A0  A1  A2  A3  S0  S1 :  X
         0   ?   ?   ?   0   0  :  0   ;
         1   ?   ?   ?   0   0  :  1   ;
         ?   0   ?   ?   1   0  :  0   ;
         ?   1   ?   ?   1   0  :  1   ;
         ?   ?   0   ?   0   1  :  0   ;
         ?   ?   1   ?   0   1  :  1   ;
         ?   ?   ?   0   1   1  :  0   ;
         ?   ?   ?   1   1   1  :  1   ;
         0   0   0   0   ?   ?  :  0   ;
         1   1   1   1   ?   ?  :  1   ;
         0   0   ?   ?   ?   0  :  0   ;
         1   1   ?   ?   ?   0  :  1   ;
         ?   ?   0   0   ?   1  :  0   ;
         ?   ?   1   1   ?   1  :  1   ;
         0   ?   0   ?   0   ?  :  0   ;
         1   ?   1   ?   0   ?  :  1   ;
         ?   0   ?   0   1   ?  :  0   ;
         ?   1   ?   1   1   ?  :  1   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_MUX_4TO2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VGND!=0
 *   UDP_OUT :=UDP_IN when VGND==0
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_pwrgood$l_pp$G (
    UDP_OUT,
    UDP_IN ,
    VGND
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VGND   ;

    table
     // UDP_IN VGND : out
          0     0   :  0   ;
          1     0   :  1   ;
          x     0   :  x   ;
          ?     1   :  x   ;
          ?     x   :  x   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_PWRGOOD_L_PP_G_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VPWR!=1 or VGND!=0
 *   UDP_OUT :=UDP_IN when VPWR==1 and VGND==0
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_pwrgood$l_pp$PG (
    UDP_OUT,
    UDP_IN ,
    VPWR   ,
    VGND
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VPWR   ;
    input  VGND   ;

    table
     // UDP_IN VPWR VGND : out
          0     1    0   :  0   ;
          1     1    0   :  1   ;
          x     1    0   :  x   ;
          ?     0    0   :  x   ;
          ?     1    1   :  x   ;
          ?     x    0   :  x   ;
          ?     1    x   :  x   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_PWRGOOD_L_PP_PG_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VPWR!=1 or VGND!=0
 *   UDP_OUT :=UDP_IN when VPWR==1 and VGND==0
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_pwrgood$l_pp$PG$S (
    UDP_OUT,
    UDP_IN ,
    VPWR   ,
    VGND   ,
    SLEEP
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VPWR   ;
    input  VGND   ;
    input  SLEEP  ;

    table
     // UDP_IN VPWR VGND SLEEP : out
          0     1    0     ?   :  0   ;
          1     1    0     0   :  1   ;
          x     1    0     0   :  x   ;
          ?     0    0     0   :  x   ;
          ?     1    1     0   :  x   ;
          ?     x    0     0   :  x   ;
          ?     1    x     0   :  x   ;
          ?     ?    0     1   :  0   ;
          ?     ?    1     1   :  x   ;
          ?     ?    x     1   :  x   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_PWRGOOD_L_PP_PG_S_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VPWR!=1
 *   UDP_OUT :=UDP_IN when VPWR==1
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_pwrgood_pp$G (
    UDP_OUT,
    UDP_IN ,
    VGND
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VGND   ;

    table
     // UDP_IN VPWR : UDP_OUT
          0     0   :    0     ;
          1     0   :    1     ;
          ?     1   :    x     ;
          ?     x   :    x     ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_PWRGOOD_PP_G_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VPWR!=1
 *   UDP_OUT :=UDP_IN when VPWR==1
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_pwrgood_pp$P (
    UDP_OUT,
    UDP_IN ,
    VPWR
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VPWR   ;

    table
     // UDP_IN VPWR : UDP_OUT
          0     1   :    0     ;
          1     1   :    1     ;
          ?     0   :    x     ;
          ?     x   :    x     ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_PWRGOOD_PP_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VPWR!=1 or VGND!=0
 *   UDP_OUT :=UDP_IN when VPWR==1 and VGND==0
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hd__udp_pwrgood_pp$PG (
    UDP_OUT,
    UDP_IN ,
    VPWR   ,
    VGND
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VPWR   ;
    input  VGND   ;

    table
     // UDP_IN VPWR VGND : out
          0     1    0   :  0   ;
          1     1    0   :  1   ;
          x     1    0   :  x   ;
          ?     0    0   :  x   ;
          ?     1    1   :  x   ;
          ?     x    0   :  x   ;
          ?     1    x   :  x   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HD__UDP_PWRGOOD_PP_PG_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2bb2o: 2-input AND, both inputs inverted, into first input, and
 *         2-input AND into 2nd input of 2-input OR.
 *
 *         X = ((!A1 & !A2) | (B1 & B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a2bb2o: 2-input AND, both inputs inverted, into first input, and
 *         2-input AND into 2nd input of 2-input OR.
 *
 *         X = ((!A1 & !A2) | (B1 & B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a2bb2o (
    X   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , B1, B2               );
    nor                                nor0        (nor0_out         , A1_N, A2_N           );
    or                                 or0         (or0_out_X        , nor0_out, and0_out   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2O_FUNCTIONAL_PP_V















































































 // FUNCTIONAL

















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2bb2o: 2-input AND, both inputs inverted, into first input, and
 *         2-input AND into 2nd input of 2-input OR.
 *
 *         X = ((!A1 & !A2) | (B1 & B2))
 *
 * Verilog wrapper for a2bb2o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2bb2o_1 (
    X   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2bb2o base (
        .X(X),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2bb2o: 2-input AND, both inputs inverted, into first input, and
 *         2-input AND into 2nd input of 2-input OR.
 *
 *         X = ((!A1 & !A2) | (B1 & B2))
 *
 * Verilog wrapper for a2bb2o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2bb2o_2 (
    X   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2bb2o base (
        .X(X),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2bb2o: 2-input AND, both inputs inverted, into first input, and
 *         2-input AND into 2nd input of 2-input OR.
 *
 *         X = ((!A1 & !A2) | (B1 & B2))
 *
 * Verilog wrapper for a2bb2o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2bb2o_4 (
    X   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2bb2o base (
        .X(X),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2bb2oi: 2-input AND, both inputs inverted, into first input, and
 *          2-input AND into 2nd input of 2-input NOR.
 *
 *          Y = !((!A1 & !A2) | (B1 & B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a2bb2oi: 2-input AND, both inputs inverted, into first input, and
 *          2-input AND into 2nd input of 2-input NOR.
 *
 *          Y = !((!A1 & !A2) | (B1 & B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a2bb2oi (
    Y   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out         ;
    wire nor1_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , B1, B2                );
    nor                                nor0        (nor0_out         , A1_N, A2_N            );
    nor                                nor1        (nor1_out_Y       , nor0_out, and0_out    );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor1_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2OI_FUNCTIONAL_PP_V















































































 // FUNCTIONAL

















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2bb2oi: 2-input AND, both inputs inverted, into first input, and
 *          2-input AND into 2nd input of 2-input NOR.
 *
 *          Y = !((!A1 & !A2) | (B1 & B2))
 *
 * Verilog wrapper for a2bb2oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2bb2oi_1 (
    Y   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2bb2oi base (
        .Y(Y),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2bb2oi: 2-input AND, both inputs inverted, into first input, and
 *          2-input AND into 2nd input of 2-input NOR.
 *
 *          Y = !((!A1 & !A2) | (B1 & B2))
 *
 * Verilog wrapper for a2bb2oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2bb2oi_2 (
    Y   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2bb2oi base (
        .Y(Y),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2bb2oi: 2-input AND, both inputs inverted, into first input, and
 *          2-input AND into 2nd input of 2-input NOR.
 *
 *          Y = !((!A1 & !A2) | (B1 & B2))
 *
 * Verilog wrapper for a2bb2oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2bb2oi_4 (
    Y   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2bb2oi base (
        .Y(Y),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2BB2OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21bo: 2-input AND into first input of 2-input OR,
 *        2nd input inverted.
 *
 *        X = ((A1 & A2) | (!B1_N))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a21bo: 2-input AND into first input of 2-input OR,
 *        2nd input inverted.
 *
 *        X = ((A1 & A2) | (!B1_N))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a21bo (
    X   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire nand1_out_X      ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out        , A2, A1                 );
    nand                               nand1       (nand1_out_X      , B1_N, nand0_out        );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, nand1_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A21BO_FUNCTIONAL_PP_V











































































 // FUNCTIONAL









































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BO_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21bo: 2-input AND into first input of 2-input OR,
 *        2nd input inverted.
 *
 *        X = ((A1 & A2) | (!B1_N))
 *
 * Verilog wrapper for a21bo with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21bo_1 (
    X   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21bo base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BO_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21bo: 2-input AND into first input of 2-input OR,
 *        2nd input inverted.
 *
 *        X = ((A1 & A2) | (!B1_N))
 *
 * Verilog wrapper for a21bo with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21bo_2 (
    X   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21bo base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BO_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21bo: 2-input AND into first input of 2-input OR,
 *        2nd input inverted.
 *
 *        X = ((A1 & A2) | (!B1_N))
 *
 * Verilog wrapper for a21bo with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21bo_4 (
    X   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21bo base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BO_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21boi: 2-input AND into first input of 2-input NOR,
 *         2nd input inverted.
 *
 *         Y = !((A1 & A2) | (!B1_N))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a21boi: 2-input AND into first input of 2-input NOR,
 *         2nd input inverted.
 *
 *         Y = !((A1 & A2) | (!B1_N))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a21boi (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire b                ;
    wire and0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (b                , B1_N                  );
    and                                and0        (and0_out         , A1, A2                );
    nor                                nor0        (nor0_out_Y       , b, and0_out           );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A21BOI_FUNCTIONAL_PP_V













































































 // FUNCTIONAL













































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BOI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21boi: 2-input AND into first input of 2-input NOR,
 *         2nd input inverted.
 *
 *         Y = !((A1 & A2) | (!B1_N))
 *
 * Verilog wrapper for a21boi with size of 0 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21boi_0 (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21boi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BOI_0_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21boi: 2-input AND into first input of 2-input NOR,
 *         2nd input inverted.
 *
 *         Y = !((A1 & A2) | (!B1_N))
 *
 * Verilog wrapper for a21boi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21boi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21boi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BOI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21boi: 2-input AND into first input of 2-input NOR,
 *         2nd input inverted.
 *
 *         Y = !((A1 & A2) | (!B1_N))
 *
 * Verilog wrapper for a21boi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21boi_2 (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21boi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BOI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21boi: 2-input AND into first input of 2-input NOR,
 *         2nd input inverted.
 *
 *         Y = !((A1 & A2) | (!B1_N))
 *
 * Verilog wrapper for a21boi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21boi_4 (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21boi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21BOI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21o: 2-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2) | B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a21o: 2-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2) | B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a21o (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A1, A2               );
    or                                 or0         (or0_out_X        , and0_out, B1         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A21O_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21o: 2-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2) | B1)
 *
 * Verilog wrapper for a21o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21o_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21o: 2-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2) | B1)
 *
 * Verilog wrapper for a21o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21o_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21o: 2-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2) | B1)
 *
 * Verilog wrapper for a21o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21o_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21oi: 2-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2) | B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a21oi: 2-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2) | B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a21oi (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A1, A2                );
    nor                                nor0        (nor0_out_Y       , B1, and0_out          );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A21OI_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21oi: 2-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2) | B1)
 *
 * Verilog wrapper for a21oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21oi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21oi: 2-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2) | B1)
 *
 * Verilog wrapper for a21oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21oi_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21oi: 2-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2) | B1)
 *
 * Verilog wrapper for a21oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a21oi_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a21oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A21OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22o: 2-input AND into both inputs of 2-input OR.
 *
 *       X = ((A1 & A2) | (B1 & B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a22o: 2-input AND into both inputs of 2-input OR.
 *
 *       X = ((A1 & A2) | (B1 & B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a22o (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire and1_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , B1, B2               );
    and                                and1        (and1_out         , A1, A2               );
    or                                 or0         (or0_out_X        , and1_out, and0_out   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A22O_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A22O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22o: 2-input AND into both inputs of 2-input OR.
 *
 *       X = ((A1 & A2) | (B1 & B2))
 *
 * Verilog wrapper for a22o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a22o_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a22o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A22O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22o: 2-input AND into both inputs of 2-input OR.
 *
 *       X = ((A1 & A2) | (B1 & B2))
 *
 * Verilog wrapper for a22o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a22o_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a22o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A22O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22o: 2-input AND into both inputs of 2-input OR.
 *
 *       X = ((A1 & A2) | (B1 & B2))
 *
 * Verilog wrapper for a22o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a22o_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a22o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A22O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22oi: 2-input AND into both inputs of 2-input NOR.
 *
 *        Y = !((A1 & A2) | (B1 & B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a22oi: 2-input AND into both inputs of 2-input NOR.
 *
 *        Y = !((A1 & A2) | (B1 & B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a22oi (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire nand1_out        ;
    wire and0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out        , A2, A1                );
    nand                               nand1       (nand1_out        , B2, B1                );
    and                                and0        (and0_out_Y       , nand0_out, nand1_out  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, and0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A22OI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A22OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22oi: 2-input AND into both inputs of 2-input NOR.
 *
 *        Y = !((A1 & A2) | (B1 & B2))
 *
 * Verilog wrapper for a22oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a22oi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a22oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A22OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22oi: 2-input AND into both inputs of 2-input NOR.
 *
 *        Y = !((A1 & A2) | (B1 & B2))
 *
 * Verilog wrapper for a22oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a22oi_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a22oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A22OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22oi: 2-input AND into both inputs of 2-input NOR.
 *
 *        Y = !((A1 & A2) | (B1 & B2))
 *
 * Verilog wrapper for a22oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a22oi_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a22oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A22OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a31o: 3-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a31o: 3-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a31o (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A3, A1, A2           );
    or                                 or0         (or0_out_X        , and0_out, B1         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A31O_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A31O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a31o: 3-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | B1)
 *
 * Verilog wrapper for a31o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a31o_1 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a31o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A31O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a31o: 3-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | B1)
 *
 * Verilog wrapper for a31o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a31o_2 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a31o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A31O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a31o: 3-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | B1)
 *
 * Verilog wrapper for a31o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a31o_4 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a31o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A31O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a31oi: 3-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a31oi: 3-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a31oi (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A3, A1, A2            );
    nor                                nor0        (nor0_out_Y       , B1, and0_out          );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A31OI_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A31OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a31oi: 3-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | B1)
 *
 * Verilog wrapper for a31oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a31oi_1 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a31oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A31OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a31oi: 3-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | B1)
 *
 * Verilog wrapper for a31oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a31oi_2 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a31oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A31OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a31oi: 3-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | B1)
 *
 * Verilog wrapper for a31oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a31oi_4 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a31oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A31OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a32o: 3-input AND into first input, and 2-input AND into
 *       2nd input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a32o: 3-input AND into first input, and 2-input AND into
 *       2nd input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a32o (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire and1_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A3, A1, A2           );
    and                                and1        (and1_out         , B1, B2               );
    or                                 or0         (or0_out_X        , and1_out, and0_out   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A32O_FUNCTIONAL_PP_V

















































































 // FUNCTIONAL





















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A32O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a32o: 3-input AND into first input, and 2-input AND into
 *       2nd input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog wrapper for a32o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a32o_1 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a32o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A32O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a32o: 3-input AND into first input, and 2-input AND into
 *       2nd input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog wrapper for a32o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a32o_2 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a32o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A32O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a32o: 3-input AND into first input, and 2-input AND into
 *       2nd input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog wrapper for a32o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a32o_4 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a32o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A32O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a32oi: 3-input AND into first input, and 2-input AND into
 *        2nd input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a32oi: 3-input AND into first input, and 2-input AND into
 *        2nd input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a32oi (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire nand1_out        ;
    wire and0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out        , A2, A1, A3            );
    nand                               nand1       (nand1_out        , B2, B1                );
    and                                and0        (and0_out_Y       , nand0_out, nand1_out  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, and0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A32OI_FUNCTIONAL_PP_V

















































































 // FUNCTIONAL





















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A32OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a32oi: 3-input AND into first input, and 2-input AND into
 *        2nd input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog wrapper for a32oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a32oi_1 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a32oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A32OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a32oi: 3-input AND into first input, and 2-input AND into
 *        2nd input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog wrapper for a32oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a32oi_2 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a32oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A32OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a32oi: 3-input AND into first input, and 2-input AND into
 *        2nd input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3) | (B1 & B2))
 *
 * Verilog wrapper for a32oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a32oi_4 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a32oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A32OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a41o: 4-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a41o: 4-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a41o (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A1, A2, A3, A4       );
    or                                 or0         (or0_out_X        , and0_out, B1         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A41O_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A41O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a41o: 4-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog wrapper for a41o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a41o_1 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a41o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A41O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a41o: 4-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog wrapper for a41o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a41o_2 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a41o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A41O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a41o: 4-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog wrapper for a41o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a41o_4 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a41o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A41O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a41oi: 4-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a41oi: 4-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a41oi (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A1, A2, A3, A4        );
    nor                                nor0        (nor0_out_Y       , B1, and0_out          );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A41OI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A41OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a41oi: 4-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog wrapper for a41oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a41oi_1 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a41oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A41OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a41oi: 4-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog wrapper for a41oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a41oi_2 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a41oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A41OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a41oi: 4-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2 & A3 & A4) | B1)
 *
 * Verilog wrapper for a41oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a41oi_4 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a41oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A41OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a211o: 2-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2) | B1 | C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a211o: 2-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2) | B1 | C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a211o (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A1, A2               );
    or                                 or0         (or0_out_X        , and0_out, C1, B1     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A211O_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A211O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a211o: 2-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2) | B1 | C1)
 *
 * Verilog wrapper for a211o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a211o_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a211o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A211O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a211o: 2-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2) | B1 | C1)
 *
 * Verilog wrapper for a211o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a211o_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a211o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A211O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a211o: 2-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2) | B1 | C1)
 *
 * Verilog wrapper for a211o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a211o_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a211o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A211O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a211oi: 2-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2) | B1 | C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a211oi: 2-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2) | B1 | C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a211oi (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A1, A2                );
    nor                                nor0        (nor0_out_Y       , and0_out, B1, C1      );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A211OI_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A211OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a211oi: 2-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2) | B1 | C1)
 *
 * Verilog wrapper for a211oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a211oi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a211oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A211OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a211oi: 2-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2) | B1 | C1)
 *
 * Verilog wrapper for a211oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a211oi_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a211oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A211OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a211oi: 2-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2) | B1 | C1)
 *
 * Verilog wrapper for a211oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a211oi_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a211oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A211OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a221o: 2-input AND into first two inputs of 3-input OR.
 *
 *        X = ((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a221o: 2-input AND into first two inputs of 3-input OR.
 *
 *        X = ((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a221o (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire and1_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , B1, B2                );
    and                                and1        (and1_out         , A1, A2                );
    or                                 or0         (or0_out_X        , and1_out, and0_out, C1);
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND );
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A221O_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL



















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A221O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a221o: 2-input AND into first two inputs of 3-input OR.
 *
 *        X = ((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog wrapper for a221o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a221o_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a221o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A221O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a221o: 2-input AND into first two inputs of 3-input OR.
 *
 *        X = ((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog wrapper for a221o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a221o_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a221o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A221O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a221o: 2-input AND into first two inputs of 3-input OR.
 *
 *        X = ((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog wrapper for a221o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a221o_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a221o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A221O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a221oi: 2-input AND into first two inputs of 3-input NOR.
 *
 *         Y = !((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a221oi: 2-input AND into first two inputs of 3-input NOR.
 *
 *         Y = !((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a221oi (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire and1_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , B1, B2                );
    and                                and1        (and1_out         , A1, A2                );
    nor                                nor0        (nor0_out_Y       , and0_out, C1, and1_out);
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A221OI_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL



















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A221OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a221oi: 2-input AND into first two inputs of 3-input NOR.
 *
 *         Y = !((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog wrapper for a221oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a221oi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a221oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A221OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a221oi: 2-input AND into first two inputs of 3-input NOR.
 *
 *         Y = !((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog wrapper for a221oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a221oi_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a221oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A221OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a221oi: 2-input AND into first two inputs of 3-input NOR.
 *
 *         Y = !((A1 & A2) | (B1 & B2) | C1)
 *
 * Verilog wrapper for a221oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a221oi_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a221oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A221OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a222oi: 2-input AND into all inputs of 3-input NOR.
 *
 *         Y = !((A1 & A2) | (B1 & B2) | (C1 & C2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a222oi: 2-input AND into all inputs of 3-input NOR.
 *
 *         Y = !((A1 & A2) | (B1 & B2) | (C1 & C2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a222oi (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    C2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  C2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire nand1_out        ;
    wire nand2_out        ;
    wire and0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out        , A2, A1                         );
    nand                               nand1       (nand1_out        , B2, B1                         );
    nand                               nand2       (nand2_out        , C2, C1                         );
    and                                and0        (and0_out_Y       , nand0_out, nand1_out, nand2_out);
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, and0_out_Y, VPWR, VGND         );
    buf                                buf0        (Y                , pwrgood_pp0_out_Y              );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A222OI_FUNCTIONAL_PP_V




















































































 // FUNCTIONAL



























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A222OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a222oi: 2-input AND into all inputs of 3-input NOR.
 *
 *         Y = !((A1 & A2) | (B1 & B2) | (C1 & C2))
 *
 * Verilog wrapper for a222oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a222oi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    C2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  C2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a222oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .C2(C2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A222OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a311o: 3-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a311o: 3-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a311o (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A3, A1, A2           );
    or                                 or0         (or0_out_X        , and0_out, C1, B1     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A311O_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A311O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a311o: 3-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog wrapper for a311o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a311o_1 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a311o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A311O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a311o: 3-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog wrapper for a311o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a311o_2 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a311o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A311O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a311o: 3-input AND into first input of 3-input OR.
 *
 *        X = ((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog wrapper for a311o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a311o_4 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a311o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A311O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a311oi: 3-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a311oi: 3-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a311oi (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A3, A1, A2            );
    nor                                nor0        (nor0_out_Y       , and0_out, B1, C1      );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A311OI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A311OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a311oi: 3-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog wrapper for a311oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a311oi_1 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a311oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A311OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a311oi: 3-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog wrapper for a311oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a311oi_2 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a311oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A311OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a311oi: 3-input AND into first input of 3-input NOR.
 *
 *         Y = !((A1 & A2 & A3) | B1 | C1)
 *
 * Verilog wrapper for a311oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a311oi_4 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a311oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A311OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111o: 2-input AND into first input of 4-input OR.
 *
 *         X = ((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a2111o: 2-input AND into first input of 4-input OR.
 *
 *         X = ((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a2111o (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A1, A2               );
    or                                 or0         (or0_out_X        , C1, B1, and0_out, D1 );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A2111O_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111o: 2-input AND into first input of 4-input OR.
 *
 *         X = ((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog wrapper for a2111o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2111o_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2111o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111o: 2-input AND into first input of 4-input OR.
 *
 *         X = ((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog wrapper for a2111o with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2111o_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2111o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111O_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111o: 2-input AND into first input of 4-input OR.
 *
 *         X = ((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog wrapper for a2111o with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2111o_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2111o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111O_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111oi: 2-input AND into first input of 4-input NOR.
 *
 *          Y = !((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a2111oi: 2-input AND into first input of 4-input NOR.
 *
 *          Y = !((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__a2111oi (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out         , A1, A2                );
    nor                                nor0        (nor0_out_Y       , B1, C1, D1, and0_out  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__A2111OI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111oi: 2-input AND into first input of 4-input NOR.
 *
 *          Y = !((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog wrapper for a2111oi with size of 0 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2111oi_0 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2111oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111OI_0_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111oi: 2-input AND into first input of 4-input NOR.
 *
 *          Y = !((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog wrapper for a2111oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2111oi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2111oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111oi: 2-input AND into first input of 4-input NOR.
 *
 *          Y = !((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog wrapper for a2111oi with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2111oi_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2111oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111OI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a2111oi: 2-input AND into first input of 4-input NOR.
 *
 *          Y = !((A1 & A2) | B1 | C1 | D1)
 *
 * Verilog wrapper for a2111oi with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__a2111oi_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__a2111oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__A2111OI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2: 2-input AND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and2: 2-input AND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__and2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out_X       , A, B                  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__AND2_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2: 2-input AND.
 *
 * Verilog wrapper for and2 with size of 0 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and2_0 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2_0_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2: 2-input AND.
 *
 * Verilog wrapper for and2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and2_1 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2: 2-input AND.
 *
 * Verilog wrapper for and2 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and2_2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2: 2-input AND.
 *
 * Verilog wrapper for and2 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and2_4 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2b: 2-input AND, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and2b: 2-input AND, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__and2b (
    X   ,
    A_N ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A_N ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , A_N                   );
    and                                and0        (and0_out_X       , not0_out, B           );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__AND2B_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2b: 2-input AND, first input inverted.
 *
 * Verilog wrapper for and2b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and2b_1 (
    X   ,
    A_N ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and2b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2b: 2-input AND, first input inverted.
 *
 * Verilog wrapper for and2b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and2b_2 (
    X   ,
    A_N ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and2b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2b: 2-input AND, first input inverted.
 *
 * Verilog wrapper for and2b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and2b_4 (
    X   ,
    A_N ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and2b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND2B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3: 3-input AND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and3: 3-input AND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__and3 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out_X       , C, A, B               );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__AND3_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3: 3-input AND.
 *
 * Verilog wrapper for and3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and3_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3: 3-input AND.
 *
 * Verilog wrapper for and3 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and3_2 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND3_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3: 3-input AND.
 *
 * Verilog wrapper for and3 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and3_4 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND3_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3b: 3-input AND, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and3b: 3-input AND, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__and3b (
    X   ,
    A_N ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , A_N                   );
    and                                and0        (and0_out_X       , C, not0_out, B        );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__AND3B_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND3B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3b: 3-input AND, first input inverted.
 *
 * Verilog wrapper for and3b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and3b_1 (
    X   ,
    A_N ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and3b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND3B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3b: 3-input AND, first input inverted.
 *
 * Verilog wrapper for and3b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and3b_2 (
    X   ,
    A_N ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and3b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND3B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3b: 3-input AND, first input inverted.
 *
 * Verilog wrapper for and3b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and3b_4 (
    X   ,
    A_N ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and3b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND3B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4: 4-input AND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and4: 4-input AND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__and4 (
    X   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    and                                and0        (and0_out_X       , A, B, C, D            );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__AND4_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4: 4-input AND.
 *
 * Verilog wrapper for and4 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4: 4-input AND.
 *
 * Verilog wrapper for and4 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4_2 (
    X   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4: 4-input AND.
 *
 * Verilog wrapper for and4 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4_4 (
    X   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4b: 4-input AND, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and4b: 4-input AND, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__and4b (
    X   ,
    A_N ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , A_N                   );
    and                                and0        (and0_out_X       , not0_out, B, C, D     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__AND4B_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4b: 4-input AND, first input inverted.
 *
 * Verilog wrapper for and4b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4b_1 (
    X   ,
    A_N ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4b: 4-input AND, first input inverted.
 *
 * Verilog wrapper for and4b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4b_2 (
    X   ,
    A_N ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4b: 4-input AND, first input inverted.
 *
 * Verilog wrapper for and4b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4b_4 (
    X   ,
    A_N ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4b base (
        .X(X),
        .A_N(A_N),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4bb: 4-input AND, first two inputs inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and4bb: 4-input AND, first two inputs inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__and4bb (
    X   ,
    A_N ,
    B_N ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A_N ;
    input  B_N ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out         ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out         , A_N, B_N              );
    and                                and0        (and0_out_X       , nor0_out, C, D        );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__AND4BB_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4BB_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4bb: 4-input AND, first two inputs inverted.
 *
 * Verilog wrapper for and4bb with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4bb_1 (
    X   ,
    A_N ,
    B_N ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B_N ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4bb base (
        .X(X),
        .A_N(A_N),
        .B_N(B_N),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4BB_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4bb: 4-input AND, first two inputs inverted.
 *
 * Verilog wrapper for and4bb with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4bb_2 (
    X   ,
    A_N ,
    B_N ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B_N ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4bb base (
        .X(X),
        .A_N(A_N),
        .B_N(B_N),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4BB_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and4bb: 4-input AND, first two inputs inverted.
 *
 * Verilog wrapper for and4bb with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__and4bb_4 (
    X   ,
    A_N ,
    B_N ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A_N ;
    input  B_N ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__and4bb base (
        .X(X),
        .A_N(A_N),
        .B_N(B_N),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__AND4BB_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * buf: Buffer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__buf (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__buf_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__buf_2 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__buf_4 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 6 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__buf_6 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_6_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__buf_8 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 12 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__buf_12 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_12_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__buf_16 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUF_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * bufbuf: Double buffer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * bufbuf: Double buffer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__bufbuf (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__BUFBUF_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUFBUF_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * bufbuf: Double buffer.
 *
 * Verilog wrapper for bufbuf with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__bufbuf_8 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__bufbuf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUFBUF_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * bufbuf: Double buffer.
 *
 * Verilog wrapper for bufbuf with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__bufbuf_16 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__bufbuf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUFBUF_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * bufinv: Buffer followed by inverter.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * bufinv: Buffer followed by inverter.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__bufinv (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out_Y       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, not0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__BUFINV_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUFINV_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * bufinv: Buffer followed by inverter.
 *
 * Verilog wrapper for bufinv with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__bufinv_8 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__bufinv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUFINV_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * bufinv: Buffer followed by inverter.
 *
 * Verilog wrapper for bufinv with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__bufinv_16 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__bufinv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__BUFINV_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkbuf: Clock tree buffer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * clkbuf: Clock tree buffer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__clkbuf (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__CLKBUF_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKBUF_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkbuf: Clock tree buffer.
 *
 * Verilog wrapper for clkbuf with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkbuf_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkbuf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKBUF_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkbuf: Clock tree buffer.
 *
 * Verilog wrapper for clkbuf with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkbuf_2 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkbuf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKBUF_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkbuf: Clock tree buffer.
 *
 * Verilog wrapper for clkbuf with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkbuf_4 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkbuf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKBUF_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkbuf: Clock tree buffer.
 *
 * Verilog wrapper for clkbuf with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkbuf_8 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkbuf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKBUF_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkbuf: Clock tree buffer.
 *
 * Verilog wrapper for clkbuf with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkbuf_16 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkbuf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKBUF_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s15: Clock Delay Buffer 4-stage 0.15um length inner stage
 *                gates.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * clkdlybuf4s15: Clock Delay Buffer 4-stage 0.15um length inner stage
 *                gates.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s15 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S15_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S15_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s15: Clock Delay Buffer 4-stage 0.15um length inner stage
 *                gates.
 *
 * Verilog wrapper for clkdlybuf4s15 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s15_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkdlybuf4s15 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S15_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s15: Clock Delay Buffer 4-stage 0.15um length inner stage
 *                gates.
 *
 * Verilog wrapper for clkdlybuf4s15 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s15_2 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkdlybuf4s15 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S15_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s18: Clock Delay Buffer 4-stage 0.18um length inner stage
 *                gates.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * clkdlybuf4s18: Clock Delay Buffer 4-stage 0.18um length inner stage
 *                gates.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s18 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S18_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S18_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s18: Clock Delay Buffer 4-stage 0.18um length inner stage
 *                gates.
 *
 * Verilog wrapper for clkdlybuf4s18 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s18_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkdlybuf4s18 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S18_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s18: Clock Delay Buffer 4-stage 0.18um length inner stage
 *                gates.
 *
 * Verilog wrapper for clkdlybuf4s18 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s18_2 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkdlybuf4s18 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S18_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s25: Clock Delay Buffer 4-stage 0.25um length inner stage
 *                gates.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * clkdlybuf4s25: Clock Delay Buffer 4-stage 0.25um length inner stage
 *                gates.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s25 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S25_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S25_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s25: Clock Delay Buffer 4-stage 0.25um length inner stage
 *                gates.
 *
 * Verilog wrapper for clkdlybuf4s25 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s25_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkdlybuf4s25 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S25_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s25: Clock Delay Buffer 4-stage 0.25um length inner stage
 *                gates.
 *
 * Verilog wrapper for clkdlybuf4s25 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s25_2 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkdlybuf4s25 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S25_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s50: Clock Delay Buffer 4-stage 0.59um length inner stage
 *                gates.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * clkdlybuf4s50: Clock Delay Buffer 4-stage 0.59um length inner stage
 *                gates.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s50 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S50_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S50_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s50: Clock Delay Buffer 4-stage 0.59um length inner stage
 *                gates.
 *
 * Verilog wrapper for clkdlybuf4s50 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s50_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkdlybuf4s50 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S50_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkdlybuf4s50: Clock Delay Buffer 4-stage 0.59um length inner stage
 *                gates.
 *
 * Verilog wrapper for clkdlybuf4s50 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkdlybuf4s50_2 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkdlybuf4s50 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKDLYBUF4S50_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinv: Clock tree inverter.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * clkinv: Clock tree inverter.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__clkinv (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out_Y       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, not0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINV_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINV_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinv: Clock tree inverter.
 *
 * Verilog wrapper for clkinv with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkinv_1 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkinv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINV_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinv: Clock tree inverter.
 *
 * Verilog wrapper for clkinv with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkinv_2 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkinv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINV_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinv: Clock tree inverter.
 *
 * Verilog wrapper for clkinv with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkinv_4 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkinv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINV_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinv: Clock tree inverter.
 *
 * Verilog wrapper for clkinv with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkinv_8 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkinv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINV_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinv: Clock tree inverter.
 *
 * Verilog wrapper for clkinv with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkinv_16 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkinv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINV_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinvlp: Lower power Clock tree inverter.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * clkinvlp: Lower power Clock tree inverter.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__clkinvlp (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out_Y       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, not0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINVLP_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINVLP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinvlp: Lower power Clock tree inverter.
 *
 * Verilog wrapper for clkinvlp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkinvlp_2 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkinvlp base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINVLP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * clkinvlp: Lower power Clock tree inverter.
 *
 * Verilog wrapper for clkinvlp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__clkinvlp_4 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__clkinvlp base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CLKINVLP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * conb: Constant value, low, high outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * conb: Constant value, low, high outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__conb (
    HI  ,
    LO  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output HI  ;
    output LO  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire pullup0_out_HI  ;
    wire pulldown0_out_LO;

    //                                Name         Output            Other arguments
    pullup                            pullup0     (pullup0_out_HI  );
    sky130_fd_sc_hd__udp_pwrgood_pp$P pwrgood_pp0 (HI              , pullup0_out_HI, VPWR  );
    pulldown                          pulldown0   (pulldown0_out_LO);
    sky130_fd_sc_hd__udp_pwrgood_pp$G pwrgood_pp1 (LO              , pulldown0_out_LO, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__CONB_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CONB_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * conb: Constant value, low, high outputs.
 *
 * Verilog wrapper for conb with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__conb_1 (
    HI  ,
    LO  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output HI  ;
    output LO  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__conb base (
        .HI(HI),
        .LO(LO),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__CONB_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__decap (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DECAP_FUNCTIONAL_PP_V



















































 // FUNCTIONAL



























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DECAP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog wrapper for decap with size of 3 units (invalid?).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__decap_3 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__decap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DECAP_3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog wrapper for decap with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__decap_4 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__decap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DECAP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog wrapper for decap with size of 6 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__decap_6 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__decap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DECAP_6_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog wrapper for decap with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__decap_8 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__decap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DECAP_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog wrapper for decap with size of 12 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__decap_12 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__decap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DECAP_12_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfbbn: Delay flop, inverted set, inverted reset, inverted clock,
 *        complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfbbn: Delay flop, inverted set, inverted reset, inverted clock,
 *        complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfbbn (
    Q      ,
    Q_N    ,
    D      ,
    CLK_N  ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  D      ;
    input  CLK_N  ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET;
    wire SET  ;
    wire CLK  ;
    wire buf_Q;

    //                                   Delay       Name  Output  Other arguments
    not                                              not0 (RESET , RESET_B                         );
    not                                              not1 (SET   , SET_B                           );
    not                                              not2 (CLK   , CLK_N                           );
    sky130_fd_sc_hd__udp_dff$NSR_pp$PG$N #1 dff0 (buf_Q , SET, RESET, CLK, D, , VPWR, VGND);
    buf                                              buf0 (Q     , buf_Q                           );
    not                                              not3 (Q_N   , buf_Q                           );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFBBN_FUNCTIONAL_PP_V





























































































 // FUNCTIONAL








































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFBBN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfbbn: Delay flop, inverted set, inverted reset, inverted clock,
 *        complementary outputs.
 *
 * Verilog wrapper for dfbbn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfbbn_1 (
    Q      ,
    Q_N    ,
    D      ,
    CLK_N  ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  D      ;
    input  CLK_N  ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfbbn base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .CLK_N(CLK_N),
        .SET_B(SET_B),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFBBN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfbbn: Delay flop, inverted set, inverted reset, inverted clock,
 *        complementary outputs.
 *
 * Verilog wrapper for dfbbn with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfbbn_2 (
    Q      ,
    Q_N    ,
    D      ,
    CLK_N  ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  D      ;
    input  CLK_N  ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfbbn base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .CLK_N(CLK_N),
        .SET_B(SET_B),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFBBN_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfbbp: Delay flop, inverted set, inverted reset,
 *        complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfbbp: Delay flop, inverted set, inverted reset,
 *        complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfbbp (
    Q      ,
    Q_N    ,
    D      ,
    CLK    ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  D      ;
    input  CLK    ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET;
    wire SET  ;
    wire buf_Q;

    //                                   Delay       Name  Output  Other arguments
    not                                              not0 (RESET , RESET_B                         );
    not                                              not1 (SET   , SET_B                           );
    sky130_fd_sc_hd__udp_dff$NSR_pp$PG$N #1 dff0 (buf_Q , SET, RESET, CLK, D, , VPWR, VGND);
    buf                                              buf0 (Q     , buf_Q                           );
    not                                              not2 (Q_N   , buf_Q                           );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFBBP_FUNCTIONAL_PP_V



























































































 // FUNCTIONAL




































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFBBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfbbp: Delay flop, inverted set, inverted reset,
 *        complementary outputs.
 *
 * Verilog wrapper for dfbbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfbbp_1 (
    Q      ,
    Q_N    ,
    D      ,
    CLK    ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  D      ;
    input  CLK    ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfbbp base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .CLK(CLK),
        .SET_B(SET_B),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFBBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrbp: Delay flop, inverted reset, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfrbp: Delay flop, inverted reset, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfrbp (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q;
    wire RESET;

    //                                  Delay       Name  Output  Other arguments
    not                                             not0 (RESET , RESET_B                    );
    sky130_fd_sc_hd__udp_dff$PR_pp$PG$N #1 dff0 (buf_Q , D, CLK, RESET, , VPWR, VGND);
    buf                                             buf0 (Q     , buf_Q                      );
    not                                             not1 (Q_N   , buf_Q                      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFRBP_FUNCTIONAL_PP_V


















































































 // FUNCTIONAL






















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrbp: Delay flop, inverted reset, complementary outputs.
 *
 * Verilog wrapper for dfrbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfrbp_1 (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfrbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrbp: Delay flop, inverted reset, complementary outputs.
 *
 * Verilog wrapper for dfrbp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfrbp_2 (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfrbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRBP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrtn: Delay flop, inverted reset, inverted clock,
 *        complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfrtn: Delay flop, inverted reset, inverted clock,
 *        complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfrtn (
    Q      ,
    CLK_N  ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  CLK_N  ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q ;
    wire RESET ;
    wire intclk;

    //                                  Delay       Name  Output  Other arguments
    not                                             not0 (RESET , RESET_B                       );
    not                                             not1 (intclk, CLK_N                         );
    sky130_fd_sc_hd__udp_dff$PR_pp$PG$N #1 dff0 (buf_Q , D, intclk, RESET, , VPWR, VGND);
    buf                                             buf0 (Q     , buf_Q                         );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFRTN_FUNCTIONAL_PP_V



















































































 // FUNCTIONAL























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRTN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrtn: Delay flop, inverted reset, inverted clock,
 *        complementary outputs.
 *
 * Verilog wrapper for dfrtn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfrtn_1 (
    Q      ,
    CLK_N  ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK_N  ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfrtn base (
        .Q(Q),
        .CLK_N(CLK_N),
        .D(D),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRTN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrtp: Delay flop, inverted reset, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfrtp: Delay flop, inverted reset, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfrtp (
    Q      ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q;
    wire RESET;

    //                                  Delay       Name  Output  Other arguments
    not                                             not0 (RESET , RESET_B                    );
    sky130_fd_sc_hd__udp_dff$PR_pp$PG$N #1 dff0 (buf_Q , D, CLK, RESET, , VPWR, VGND);
    buf                                             buf0 (Q     , buf_Q                      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFRTP_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL

















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrtp: Delay flop, inverted reset, single output.
 *
 * Verilog wrapper for dfrtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfrtp_1 (
    Q      ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfrtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrtp: Delay flop, inverted reset, single output.
 *
 * Verilog wrapper for dfrtp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfrtp_2 (
    Q      ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfrtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRTP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrtp: Delay flop, inverted reset, single output.
 *
 * Verilog wrapper for dfrtp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfrtp_4 (
    Q      ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dfrtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFRTP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfsbp: Delay flop, inverted set, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfsbp: Delay flop, inverted set, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfsbp (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf_Q;
    wire SET  ;

    //                                  Delay       Name  Output  Other arguments
    not                                             not0 (SET   , SET_B                    );
    sky130_fd_sc_hd__udp_dff$PS_pp$PG$N #1 dff0 (buf_Q , D, CLK, SET, , VPWR, VGND);
    buf                                             buf0 (Q     , buf_Q                    );
    not                                             not1 (Q_N   , buf_Q                    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFSBP_FUNCTIONAL_PP_V



















































































 // FUNCTIONAL























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFSBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfsbp: Delay flop, inverted set, complementary outputs.
 *
 * Verilog wrapper for dfsbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfsbp_1 (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__dfsbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFSBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfsbp: Delay flop, inverted set, complementary outputs.
 *
 * Verilog wrapper for dfsbp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfsbp_2 (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__dfsbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFSBP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfstp: Delay flop, inverted set, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfstp: Delay flop, inverted set, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfstp (
    Q    ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf_Q;
    wire SET  ;

    //                                  Delay       Name  Output  Other arguments
    not                                             not0 (SET   , SET_B                    );
    sky130_fd_sc_hd__udp_dff$PS_pp$PG$N #1 dff0 (buf_Q , D, CLK, SET, , VPWR, VGND);
    buf                                             buf0 (Q     , buf_Q                    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFSTP_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL

















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFSTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfstp: Delay flop, inverted set, single output.
 *
 * Verilog wrapper for dfstp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfstp_1 (
    Q    ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__dfstp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFSTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfstp: Delay flop, inverted set, single output.
 *
 * Verilog wrapper for dfstp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfstp_2 (
    Q    ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__dfstp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFSTP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfstp: Delay flop, inverted set, single output.
 *
 * Verilog wrapper for dfstp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfstp_4 (
    Q    ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__dfstp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFSTP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxbp: Delay flop, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfxbp: Delay flop, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfxbp (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q;

    //                                 Delay       Name  Output  Other arguments
    sky130_fd_sc_hd__udp_dff$P_pp$PG$N #1 dff0 (buf_Q , D, CLK, , VPWR, VGND);
    buf                                            buf0 (Q     , buf_Q               );
    not                                            not0 (Q_N   , buf_Q               );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFXBP_FUNCTIONAL_PP_V










































































 // FUNCTIONAL










































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFXBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxbp: Delay flop, complementary outputs.
 *
 * Verilog wrapper for dfxbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfxbp_1 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFXBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxbp: Delay flop, complementary outputs.
 *
 * Verilog wrapper for dfxbp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfxbp_2 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFXBP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxtp: Delay flop, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfxtp: Delay flop, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dfxtp (
    Q   ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q;

    //                                 Delay       Name  Output  Other arguments
    sky130_fd_sc_hd__udp_dff$P_pp$PG$N #1 dff0 (buf_Q , D, CLK, , VPWR, VGND);
    buf                                            buf0 (Q     , buf_Q               );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DFXTP_FUNCTIONAL_PP_V







































































 // FUNCTIONAL




































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxtp: Delay flop, single output.
 *
 * Verilog wrapper for dfxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfxtp_1 (
    Q   ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxtp: Delay flop, single output.
 *
 * Verilog wrapper for dfxtp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfxtp_2 (
    Q   ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFXTP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxtp: Delay flop, single output.
 *
 * Verilog wrapper for dfxtp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dfxtp_4 (
    Q   ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DFXTP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * diode: Antenna tie-down diode.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * diode: Antenna tie-down diode.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__diode (
    DIODE,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    input DIODE;
    input VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DIODE_FUNCTIONAL_PP_V





















































 // FUNCTIONAL





































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DIODE_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * diode: Antenna tie-down diode.
 *
 * Verilog wrapper for diode with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__diode_2 (
    DIODE,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    input DIODE;
    input VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__diode base (
        .DIODE(DIODE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/
























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DIODE_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlclkp: Clock gate.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlclkp: Clock gate.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlclkp (
    GCLK,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output GCLK;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire m0  ;
    wire clkn;

    //                                    Name     Output  Other arguments
    not                                   not0    (clkn  , CLK                     );
    sky130_fd_sc_hd__udp_dlatch$P_pp$PG$N dlatch0 (m0    , GATE, clkn, , VPWR, VGND);
    and                                   and0    (GCLK  , m0, CLK                 );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLCLKP_FUNCTIONAL_PP_V









































































 // FUNCTIONAL








































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLCLKP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlclkp: Clock gate.
 *
 * Verilog wrapper for dlclkp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlclkp_1 (
    GCLK,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output GCLK;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlclkp base (
        .GCLK(GCLK),
        .GATE(GATE),
        .CLK(CLK),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLCLKP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlclkp: Clock gate.
 *
 * Verilog wrapper for dlclkp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlclkp_2 (
    GCLK,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output GCLK;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlclkp base (
        .GCLK(GCLK),
        .GATE(GATE),
        .CLK(CLK),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLCLKP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlclkp: Clock gate.
 *
 * Verilog wrapper for dlclkp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlclkp_4 (
    GCLK,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output GCLK;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlclkp base (
        .GCLK(GCLK),
        .GATE(GATE),
        .CLK(CLK),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLCLKP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrbn: Delay latch, inverted reset, inverted enable,
 *        complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlrbn: Delay latch, inverted reset, inverted enable,
 *        complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlrbn (
    Q      ,
    Q_N    ,
    RESET_B,
    D      ,
    GATE_N ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  RESET_B;
    input  D      ;
    input  GATE_N ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET  ;
    wire intgate;
    wire buf_Q  ;

    //                                     Delay       Name     Output   Other arguments
    not                                                not0    (RESET  , RESET_B                        );
    not                                                not1    (intgate, GATE_N                         );
    sky130_fd_sc_hd__udp_dlatch$PR_pp$PG$N #1 dlatch0 (buf_Q  , D, intgate, RESET, , VPWR, VGND);
    buf                                                buf0    (Q      , buf_Q                          );
    not                                                not2    (Q_N    , buf_Q                          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLRBN_FUNCTIONAL_PP_V























































































 // FUNCTIONAL






























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRBN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrbn: Delay latch, inverted reset, inverted enable,
 *        complementary outputs.
 *
 * Verilog wrapper for dlrbn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrbn_1 (
    Q      ,
    Q_N    ,
    RESET_B,
    D      ,
    GATE_N ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  RESET_B;
    input  D      ;
    input  GATE_N ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrbn base (
        .Q(Q),
        .Q_N(Q_N),
        .RESET_B(RESET_B),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRBN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrbn: Delay latch, inverted reset, inverted enable,
 *        complementary outputs.
 *
 * Verilog wrapper for dlrbn with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrbn_2 (
    Q      ,
    Q_N    ,
    RESET_B,
    D      ,
    GATE_N ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  RESET_B;
    input  D      ;
    input  GATE_N ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrbn base (
        .Q(Q),
        .Q_N(Q_N),
        .RESET_B(RESET_B),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRBN_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrbp: Delay latch, inverted reset, non-inverted enable,
 *        complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlrbp: Delay latch, inverted reset, non-inverted enable,
 *        complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlrbp (
    Q      ,
    Q_N    ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET;
    wire buf_Q;

    //                                     Delay       Name     Output  Other arguments
    not                                                not0    (RESET , RESET_B                     );
    sky130_fd_sc_hd__udp_dlatch$PR_pp$PG$N #1 dlatch0 (buf_Q , D, GATE, RESET, , VPWR, VGND);
    buf                                                buf0    (Q     , buf_Q                       );
    not                                                not1    (Q_N   , buf_Q                       );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLRBP_FUNCTIONAL_PP_V





















































































 // FUNCTIONAL


























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrbp: Delay latch, inverted reset, non-inverted enable,
 *        complementary outputs.
 *
 * Verilog wrapper for dlrbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrbp_1 (
    Q      ,
    Q_N    ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrbp base (
        .Q(Q),
        .Q_N(Q_N),
        .RESET_B(RESET_B),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrbp: Delay latch, inverted reset, non-inverted enable,
 *        complementary outputs.
 *
 * Verilog wrapper for dlrbp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrbp_2 (
    Q      ,
    Q_N    ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrbp base (
        .Q(Q),
        .Q_N(Q_N),
        .RESET_B(RESET_B),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRBP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtn: Delay latch, inverted reset, inverted enable, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlrtn: Delay latch, inverted reset, inverted enable, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlrtn (
    Q      ,
    RESET_B,
    D      ,
    GATE_N ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE_N ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET  ;
    wire intgate;
    wire buf_Q  ;

    //                                     Delay       Name     Output   Other arguments
    not                                                not0    (RESET  , RESET_B                        );
    not                                                not1    (intgate, GATE_N                         );
    sky130_fd_sc_hd__udp_dlatch$PR_pp$PG$N #1 dlatch0 (buf_Q  , D, intgate, RESET, , VPWR, VGND);
    buf                                                buf0    (Q      , buf_Q                          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTN_FUNCTIONAL_PP_V



















































































 // FUNCTIONAL






















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtn: Delay latch, inverted reset, inverted enable, single output.
 *
 * Verilog wrapper for dlrtn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrtn_1 (
    Q      ,
    RESET_B,
    D      ,
    GATE_N ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE_N ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrtn base (
        .Q(Q),
        .RESET_B(RESET_B),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtn: Delay latch, inverted reset, inverted enable, single output.
 *
 * Verilog wrapper for dlrtn with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrtn_2 (
    Q      ,
    RESET_B,
    D      ,
    GATE_N ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE_N ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrtn base (
        .Q(Q),
        .RESET_B(RESET_B),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTN_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtn: Delay latch, inverted reset, inverted enable, single output.
 *
 * Verilog wrapper for dlrtn with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrtn_4 (
    Q      ,
    RESET_B,
    D      ,
    GATE_N ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE_N ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrtn base (
        .Q(Q),
        .RESET_B(RESET_B),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTN_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtp: Delay latch, inverted reset, non-inverted enable,
 *        single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlrtp: Delay latch, inverted reset, non-inverted enable,
 *        single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlrtp (
    Q      ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET;
    wire buf_Q;

    //                                     Delay       Name     Output  Other arguments
    not                                                not0    (RESET , RESET_B                     );
    sky130_fd_sc_hd__udp_dlatch$PR_pp$PG$N #1 dlatch0 (buf_Q , D, GATE, RESET, , VPWR, VGND);
    buf                                                buf0    (Q     , buf_Q                       );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTP_FUNCTIONAL_PP_V


















































































 // FUNCTIONAL




















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtp: Delay latch, inverted reset, non-inverted enable,
 *        single output.
 *
 * Verilog wrapper for dlrtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrtp_1 (
    Q      ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrtp base (
        .Q(Q),
        .RESET_B(RESET_B),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtp: Delay latch, inverted reset, non-inverted enable,
 *        single output.
 *
 * Verilog wrapper for dlrtp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrtp_2 (
    Q      ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrtp base (
        .Q(Q),
        .RESET_B(RESET_B),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtp: Delay latch, inverted reset, non-inverted enable,
 *        single output.
 *
 * Verilog wrapper for dlrtp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlrtp_4 (
    Q      ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__dlrtp base (
        .Q(Q),
        .RESET_B(RESET_B),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLRTP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxbn: Delay latch, inverted enable, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlxbn: Delay latch, inverted enable, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlxbn (
    Q     ,
    Q_N   ,
    D     ,
    GATE_N,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    // Module ports
    output Q     ;
    output Q_N   ;
    input  D     ;
    input  GATE_N;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;

    // Local signals
    wire GATE ;
    wire buf_Q;

    //                                    Delay       Name     Output  Other arguments
    not                                               not0    (GATE  , GATE_N               );
    sky130_fd_sc_hd__udp_dlatch$P_pp$PG$N #1 dlatch0 (buf_Q , D, GATE, , VPWR, VGND);
    buf                                               buf0    (Q     , buf_Q                );
    not                                               not1    (Q_N   , buf_Q                );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLXBN_FUNCTIONAL_PP_V












































































 // FUNCTIONAL














































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXBN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxbn: Delay latch, inverted enable, complementary outputs.
 *
 * Verilog wrapper for dlxbn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlxbn_1 (
    Q     ,
    Q_N   ,
    D     ,
    GATE_N,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    output Q     ;
    output Q_N   ;
    input  D     ;
    input  GATE_N;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;
    sky130_fd_sc_hd__dlxbn base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXBN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxbn: Delay latch, inverted enable, complementary outputs.
 *
 * Verilog wrapper for dlxbn with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlxbn_2 (
    Q     ,
    Q_N   ,
    D     ,
    GATE_N,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    output Q     ;
    output Q_N   ;
    input  D     ;
    input  GATE_N;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;
    sky130_fd_sc_hd__dlxbn base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXBN_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxbp: Delay latch, non-inverted enable, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlxbp: Delay latch, non-inverted enable, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlxbp (
    Q   ,
    Q_N ,
    D   ,
    GATE,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    output Q_N ;
    input  D   ;
    input  GATE;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q;

    //                                    Delay       Name     Output  Other arguments
    sky130_fd_sc_hd__udp_dlatch$P_pp$PG$N #1 dlatch0 (buf_Q , D, GATE, , VPWR, VGND);
    buf                                               buf0    (Q     , buf_Q                );
    not                                               not0    (Q_N   , buf_Q                );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLXBP_FUNCTIONAL_PP_V










































































 // FUNCTIONAL










































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxbp: Delay latch, non-inverted enable, complementary outputs.
 *
 * Verilog wrapper for dlxbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlxbp_1 (
    Q   ,
    Q_N ,
    D   ,
    GATE,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  D   ;
    input  GATE;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxtn: Delay latch, inverted enable, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlxtn: Delay latch, inverted enable, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlxtn (
    Q     ,
    D     ,
    GATE_N,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    // Module ports
    output Q     ;
    input  D     ;
    input  GATE_N;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;

    // Local signals
    wire GATE ;
    wire buf_Q;

    //                                    Name     Output  Other arguments
    not                                   not0    (GATE  , GATE_N               );
    sky130_fd_sc_hd__udp_dlatch$P_pp$PG$N dlatch0 (buf_Q , D, GATE, , VPWR, VGND);
    buf                                   buf0    (Q     , buf_Q                );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLXTN_FUNCTIONAL_PP_V









































































 // FUNCTIONAL








































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXTN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxtn: Delay latch, inverted enable, single output.
 *
 * Verilog wrapper for dlxtn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlxtn_1 (
    Q     ,
    D     ,
    GATE_N,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    output Q     ;
    input  D     ;
    input  GATE_N;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;
    sky130_fd_sc_hd__dlxtn base (
        .Q(Q),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXTN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxtn: Delay latch, inverted enable, single output.
 *
 * Verilog wrapper for dlxtn with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlxtn_2 (
    Q     ,
    D     ,
    GATE_N,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    output Q     ;
    input  D     ;
    input  GATE_N;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;
    sky130_fd_sc_hd__dlxtn base (
        .Q(Q),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXTN_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxtn: Delay latch, inverted enable, single output.
 *
 * Verilog wrapper for dlxtn with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlxtn_4 (
    Q     ,
    D     ,
    GATE_N,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    output Q     ;
    input  D     ;
    input  GATE_N;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;
    sky130_fd_sc_hd__dlxtn base (
        .Q(Q),
        .D(D),
        .GATE_N(GATE_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXTN_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxtp: Delay latch, non-inverted enable, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlxtp: Delay latch, non-inverted enable, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlxtp (
    Q   ,
    D   ,
    GATE,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  D   ;
    input  GATE;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q;

    //                                    Name     Output  Other arguments
    sky130_fd_sc_hd__udp_dlatch$P_pp$PG$N dlatch0 (buf_Q , D, GATE, , VPWR, VGND);
    buf                                   buf0    (Q     , buf_Q                );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLXTP_FUNCTIONAL_PP_V







































































 // FUNCTIONAL




































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxtp: Delay latch, non-inverted enable, single output.
 *
 * Verilog wrapper for dlxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlxtp_1 (
    Q   ,
    D   ,
    GATE,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  D   ;
    input  GATE;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlxtp base (
        .Q(Q),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlygate4sd1: Delay Buffer 4-stage 0.15um length inner stage gates.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlygate4sd1: Delay Buffer 4-stage 0.15um length inner stage gates.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlygate4sd1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD1_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlygate4sd1: Delay Buffer 4-stage 0.15um length inner stage gates.
 *
 * Verilog wrapper for dlygate4sd1 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlygate4sd1_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlygate4sd1 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD1_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlygate4sd2: Delay Buffer 4-stage 0.18um length inner stage gates.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlygate4sd2: Delay Buffer 4-stage 0.18um length inner stage gates.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlygate4sd2 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD2_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlygate4sd2: Delay Buffer 4-stage 0.18um length inner stage gates.
 *
 * Verilog wrapper for dlygate4sd2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlygate4sd2_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlygate4sd2 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlygate4sd3: Delay Buffer 4-stage 0.50um length inner stage gates.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlygate4sd3: Delay Buffer 4-stage 0.50um length inner stage gates.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlygate4sd3 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD3_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlygate4sd3: Delay Buffer 4-stage 0.50um length inner stage gates.
 *
 * Verilog wrapper for dlygate4sd3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlygate4sd3_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlygate4sd3 base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYGATE4SD3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlymetal6s2s: 6-inverter delay with output from 2nd stage on
 *               horizontal route.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlymetal6s2s: 6-inverter delay with output from 2nd stage on
 *               horizontal route.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlymetal6s2s (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S2S_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S2S_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlymetal6s2s: 6-inverter delay with output from 2nd stage on
 *               horizontal route.
 *
 * Verilog wrapper for dlymetal6s2s with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlymetal6s2s_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlymetal6s2s base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S2S_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlymetal6s4s: 6-inverter delay with output from 4th inverter on
 *               horizontal route.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlymetal6s4s: 6-inverter delay with output from 4th inverter on
 *               horizontal route.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlymetal6s4s (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S4S_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S4S_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlymetal6s4s: 6-inverter delay with output from 4th inverter on
 *               horizontal route.
 *
 * Verilog wrapper for dlymetal6s4s with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlymetal6s4s_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlymetal6s4s base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S4S_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlymetal6s6s: 6-inverter delay with output from 6th inverter on
 *               horizontal route.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlymetal6s6s: 6-inverter delay with output from 6th inverter on
 *               horizontal route.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__dlymetal6s6s (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S6S_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S6S_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlymetal6s6s: 6-inverter delay with output from 6th inverter on
 *               horizontal route.
 *
 * Verilog wrapper for dlymetal6s6s with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__dlymetal6s6s_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__dlymetal6s6s base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__DLYMETAL6S6S_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ebufn: Tri-state buffer, negative enable.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * ebufn: Tri-state buffer, negative enable.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__ebufn (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire pwrgood_pp0_out_A  ;
    wire pwrgood_pp1_out_teb;

    //                                 Name         Output               Other arguments
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A  , A, VPWR, VGND                         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_teb, TE_B, VPWR, VGND                      );
    bufif0                             bufif00     (Z                  , pwrgood_pp0_out_A, pwrgood_pp1_out_teb);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__EBUFN_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EBUFN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ebufn: Tri-state buffer, negative enable.
 *
 * Verilog wrapper for ebufn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__ebufn_1 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__ebufn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EBUFN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ebufn: Tri-state buffer, negative enable.
 *
 * Verilog wrapper for ebufn with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__ebufn_2 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__ebufn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EBUFN_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ebufn: Tri-state buffer, negative enable.
 *
 * Verilog wrapper for ebufn with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__ebufn_4 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__ebufn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EBUFN_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ebufn: Tri-state buffer, negative enable.
 *
 * Verilog wrapper for ebufn with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__ebufn_8 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__ebufn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EBUFN_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * edfxbp: Delay flop with loopback enable, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * edfxbp: Delay flop with loopback enable, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__edfxbp (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    DE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q  ;
    wire mux_out;

    //                                 Delay       Name       Output   Other arguments
    sky130_fd_sc_hd__udp_mux_2to1                  mux_2to10 (mux_out, buf_Q, D, DE              );
    sky130_fd_sc_hd__udp_dff$P_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, , VPWR, VGND);
    buf                                            buf0      (Q      , buf_Q                     );
    not                                            not0      (Q_N    , buf_Q                     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__EDFXBP_FUNCTIONAL_PP_V


















































































 // FUNCTIONAL























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EDFXBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * edfxbp: Delay flop with loopback enable, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog wrapper for edfxbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__edfxbp_1 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    DE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__edfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .DE(DE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EDFXBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * edfxtp: Delay flop with loopback enable, non-inverted clock,
 *         single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * edfxtp: Delay flop with loopback enable, non-inverted clock,
 *         single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__edfxtp (
    Q   ,
    CLK ,
    D   ,
    DE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q  ;
    wire mux_out;

    //                                 Delay       Name       Output   Other arguments
    sky130_fd_sc_hd__udp_mux_2to1                  mux_2to10 (mux_out, buf_Q, D, DE              );
    sky130_fd_sc_hd__udp_dff$P_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, , VPWR, VGND);
    buf                                            buf0      (Q      , buf_Q                     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__EDFXTP_FUNCTIONAL_PP_V















































































 // FUNCTIONAL

















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EDFXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * edfxtp: Delay flop with loopback enable, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for edfxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__edfxtp_1 (
    Q   ,
    CLK ,
    D   ,
    DE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__edfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .DE(DE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EDFXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__einvn (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire pwrgood_pp0_out_A  ;
    wire pwrgood_pp1_out_teb;

    //                                 Name         Output               Other arguments
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A  , A, VPWR, VGND                         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_teb, TE_B, VPWR, VGND                      );
    notif0                             notif00     (Z                  , pwrgood_pp0_out_A, pwrgood_pp1_out_teb);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__EINVN_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog wrapper for einvn with size of 0 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvn_0 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVN_0_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog wrapper for einvn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvn_1 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog wrapper for einvn with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvn_2 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVN_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog wrapper for einvn with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvn_4 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVN_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog wrapper for einvn with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvn_8 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVN_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__einvp (
    Z   ,
    A   ,
    TE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Z   ;
    input  A   ;
    input  TE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire pwrgood_pp0_out_A ;
    wire pwrgood_pp1_out_TE;

    //                                 Name         Output              Other arguments
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A , A, VPWR, VGND                        );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_TE, TE, VPWR, VGND                       );
    notif1                             notif10     (Z                 , pwrgood_pp0_out_A, pwrgood_pp1_out_TE);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__EINVP_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog wrapper for einvp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvp_1 (
    Z   ,
    A   ,
    TE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvp base (
        .Z(Z),
        .A(A),
        .TE(TE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog wrapper for einvp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvp_2 (
    Z   ,
    A   ,
    TE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvp base (
        .Z(Z),
        .A(A),
        .TE(TE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog wrapper for einvp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvp_4 (
    Z   ,
    A   ,
    TE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvp base (
        .Z(Z),
        .A(A),
        .TE(TE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog wrapper for einvp with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__einvp_8 (
    Z   ,
    A   ,
    TE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__einvp base (
        .Z(Z),
        .A(A),
        .TE(TE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__EINVP_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fa: Full adder.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * fa: Full adder.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__fa (
    COUT,
    SUM ,
    A   ,
    B   ,
    CIN ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  CIN ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out             ;
    wire and0_out            ;
    wire and1_out            ;
    wire and2_out            ;
    wire nor0_out            ;
    wire nor1_out            ;
    wire or1_out_COUT        ;
    wire pwrgood_pp0_out_COUT;
    wire or2_out_SUM         ;
    wire pwrgood_pp1_out_SUM ;

    //                                 Name         Output                Other arguments
    or                                 or0         (or0_out             , CIN, B                  );
    and                                and0        (and0_out            , or0_out, A              );
    and                                and1        (and1_out            , B, CIN                  );
    or                                 or1         (or1_out_COUT        , and1_out, and0_out      );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_COUT, or1_out_COUT, VPWR, VGND);
    buf                                buf0        (COUT                , pwrgood_pp0_out_COUT    );
    and                                and2        (and2_out            , CIN, A, B               );
    nor                                nor0        (nor0_out            , A, or0_out              );
    nor                                nor1        (nor1_out            , nor0_out, COUT          );
    or                                 or2         (or2_out_SUM         , nor1_out, and2_out      );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_SUM , or2_out_SUM, VPWR, VGND );
    buf                                buf1        (SUM                 , pwrgood_pp1_out_SUM     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__FA_FUNCTIONAL_PP_V

























































































 // FUNCTIONAL

































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FA_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fa: Full adder.
 *
 * Verilog wrapper for fa with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fa_1 (
    COUT,
    SUM ,
    A   ,
    B   ,
    CIN ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  CIN ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__fa base (
        .COUT(COUT),
        .SUM(SUM),
        .A(A),
        .B(B),
        .CIN(CIN),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FA_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fa: Full adder.
 *
 * Verilog wrapper for fa with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fa_2 (
    COUT,
    SUM ,
    A   ,
    B   ,
    CIN ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  CIN ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__fa base (
        .COUT(COUT),
        .SUM(SUM),
        .A(A),
        .B(B),
        .CIN(CIN),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FA_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fa: Full adder.
 *
 * Verilog wrapper for fa with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fa_4 (
    COUT,
    SUM ,
    A   ,
    B   ,
    CIN ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  CIN ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__fa base (
        .COUT(COUT),
        .SUM(SUM),
        .A(A),
        .B(B),
        .CIN(CIN),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FA_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fah: Full adder.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * fah: Full adder.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__fah (
    COUT,
    SUM ,
    A   ,
    B   ,
    CI  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  CI  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire xor0_out_SUM        ;
    wire pwrgood_pp0_out_SUM ;
    wire a_b                 ;
    wire a_ci                ;
    wire b_ci                ;
    wire or0_out_COUT        ;
    wire pwrgood_pp1_out_COUT;

    //                                 Name         Output                Other arguments
    xor                                xor0        (xor0_out_SUM        , A, B, CI                );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_SUM , xor0_out_SUM, VPWR, VGND);
    buf                                buf0        (SUM                 , pwrgood_pp0_out_SUM     );
    and                                and0        (a_b                 , A, B                    );
    and                                and1        (a_ci                , A, CI                   );
    and                                and2        (b_ci                , B, CI                   );
    or                                 or0         (or0_out_COUT        , a_b, a_ci, b_ci         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_COUT, or0_out_COUT, VPWR, VGND);
    buf                                buf1        (COUT                , pwrgood_pp1_out_COUT    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__FAH_FUNCTIONAL_PP_V



















































































 // FUNCTIONAL





















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FAH_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fah: Full adder.
 *
 * Verilog wrapper for fah with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fah_1 (
    COUT,
    SUM ,
    A   ,
    B   ,
    CI  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  CI  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__fah base (
        .COUT(COUT),
        .SUM(SUM),
        .A(A),
        .B(B),
        .CI(CI),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FAH_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fahcin: Full adder, inverted carry in.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * fahcin: Full adder, inverted carry in.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__fahcin (
    COUT,
    SUM ,
    A   ,
    B   ,
    CIN ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  CIN ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire ci                  ;
    wire xor0_out_SUM        ;
    wire pwrgood_pp0_out_SUM ;
    wire a_b                 ;
    wire a_ci                ;
    wire b_ci                ;
    wire or0_out_COUT        ;
    wire pwrgood_pp1_out_COUT;

    //                                 Name         Output                Other arguments
    not                                not0        (ci                  , CIN                     );
    xor                                xor0        (xor0_out_SUM        , A, B, ci                );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_SUM , xor0_out_SUM, VPWR, VGND);
    buf                                buf0        (SUM                 , pwrgood_pp0_out_SUM     );
    and                                and0        (a_b                 , A, B                    );
    and                                and1        (a_ci                , A, ci                   );
    and                                and2        (b_ci                , B, ci                   );
    or                                 or0         (or0_out_COUT        , a_b, a_ci, b_ci         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_COUT, or0_out_COUT, VPWR, VGND);
    buf                                buf1        (COUT                , pwrgood_pp1_out_COUT    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__FAHCIN_FUNCTIONAL_PP_V





















































































 // FUNCTIONAL

























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FAHCIN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fahcin: Full adder, inverted carry in.
 *
 * Verilog wrapper for fahcin with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fahcin_1 (
    COUT,
    SUM ,
    A   ,
    B   ,
    CIN ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  CIN ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__fahcin base (
        .COUT(COUT),
        .SUM(SUM),
        .A(A),
        .B(B),
        .CIN(CIN),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FAHCIN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fahcon: Full adder, inverted carry in, inverted carry out.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * fahcon: Full adder, inverted carry in, inverted carry out.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__fahcon (
    COUT_N,
    SUM   ,
    A     ,
    B     ,
    CI    ,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    // Module ports
    output COUT_N;
    output SUM   ;
    input  A     ;
    input  B     ;
    input  CI    ;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;

    // Local signals
    wire xor0_out_SUM         ;
    wire pwrgood_pp0_out_SUM  ;
    wire a_b                  ;
    wire a_ci                 ;
    wire b_ci                 ;
    wire or0_out_coutn        ;
    wire pwrgood_pp1_out_coutn;

    //                                 Name         Output                 Other arguments
    xor                                xor0        (xor0_out_SUM         , A, B, CI                 );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_SUM  , xor0_out_SUM, VPWR, VGND );
    buf                                buf0        (SUM                  , pwrgood_pp0_out_SUM      );
    nor                                nor0        (a_b                  , A, B                     );
    nor                                nor1        (a_ci                 , A, CI                    );
    nor                                nor2        (b_ci                 , B, CI                    );
    or                                 or0         (or0_out_coutn        , a_b, a_ci, b_ci          );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_coutn, or0_out_coutn, VPWR, VGND);
    buf                                buf1        (COUT_N               , pwrgood_pp1_out_coutn    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__FAHCON_FUNCTIONAL_PP_V



















































































 // FUNCTIONAL





















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FAHCON_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fahcon: Full adder, inverted carry in, inverted carry out.
 *
 * Verilog wrapper for fahcon with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fahcon_1 (
    COUT_N,
    SUM   ,
    A     ,
    B     ,
    CI    ,
    VPWR  ,
    VGND  ,
    VPB   ,
    VNB
);

    output COUT_N;
    output SUM   ;
    input  A     ;
    input  B     ;
    input  CI    ;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    input  VNB   ;
    sky130_fd_sc_hd__fahcon base (
        .COUT_N(COUT_N),
        .SUM(SUM),
        .A(A),
        .B(B),
        .CI(CI),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FAHCON_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * fill: Fill cell.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__fill (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__FILL_FUNCTIONAL_PP_V



















































 // FUNCTIONAL

































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FILL_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fill_1 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FILL_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fill_2 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FILL_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fill_4 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FILL_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__fill_8 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__FILL_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ha: Half adder.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * ha: Half adder.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__ha (
    COUT,
    SUM ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out_COUT       ;
    wire pwrgood_pp0_out_COUT;
    wire xor0_out_SUM        ;
    wire pwrgood_pp1_out_SUM ;

    //                                 Name         Output                Other arguments
    and                                and0        (and0_out_COUT       , A, B                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_COUT, and0_out_COUT, VPWR, VGND);
    buf                                buf0        (COUT                , pwrgood_pp0_out_COUT     );
    xor                                xor0        (xor0_out_SUM        , B, A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_SUM , xor0_out_SUM, VPWR, VGND );
    buf                                buf1        (SUM                 , pwrgood_pp1_out_SUM      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__HA_FUNCTIONAL_PP_V











































































 // FUNCTIONAL





































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__HA_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ha: Half adder.
 *
 * Verilog wrapper for ha with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__ha_1 (
    COUT,
    SUM ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__ha base (
        .COUT(COUT),
        .SUM(SUM),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__HA_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ha: Half adder.
 *
 * Verilog wrapper for ha with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__ha_2 (
    COUT,
    SUM ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__ha base (
        .COUT(COUT),
        .SUM(SUM),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__HA_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * ha: Half adder.
 *
 * Verilog wrapper for ha with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__ha_4 (
    COUT,
    SUM ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output COUT;
    output SUM ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__ha base (
        .COUT(COUT),
        .SUM(SUM),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__HA_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * inv: Inverter.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__inv (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out_Y       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, not0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__INV_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__INV_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__inv_1 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__INV_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__inv_2 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__INV_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__inv_4 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__INV_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 6 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__inv_6 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__INV_6_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__inv_8 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__INV_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 12 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__inv_12 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__INV_12_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__inv_16 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__INV_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_bleeder: Current bleeder (weak pulldown to ground).
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/




`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__lpflow_bleeder (
    SHORT,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    input SHORT;
    inout VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;

endmodule
`endcelldefine

`default_nettype wire
	// SKY130_FD_SC_HD__LPFLOW_BLEEDER_FUNCTIONAL_PP_V


















































 // FUNCTIONAL















































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_BLEEDER_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_bleeder: Current bleeder (weak pulldown to ground).
 *
 * Verilog wrapper for lpflow_bleeder with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_bleeder_1 (
    SHORT,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    input SHORT;
    inout VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__lpflow_bleeder base (
        .SHORT(SHORT),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/
























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_BLEEDER_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkbufkapwr: Clock tree buffer on keep-alive power rail.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_clkbufkapwr: Clock tree buffer on keep-alive power rail.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_clkbufkapwr (
    X    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf0_out_X    ;
    wire pwrgood0_out_X;

    //                                   Name      Output          Other arguments
    buf                                  buf0     (buf0_out_X    , A                      );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (pwrgood0_out_X, buf0_out_X, KAPWR, VGND);
    buf                                  buf1     (X             , pwrgood0_out_X         );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_FUNCTIONAL_PP_V




































































 // FUNCTIONAL
























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkbufkapwr: Clock tree buffer on keep-alive power rail.
 *
 * Verilog wrapper for lpflow_clkbufkapwr with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkbufkapwr_1 (
    X    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkbufkapwr base (
        .X(X),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkbufkapwr: Clock tree buffer on keep-alive power rail.
 *
 * Verilog wrapper for lpflow_clkbufkapwr with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkbufkapwr_2 (
    X    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkbufkapwr base (
        .X(X),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkbufkapwr: Clock tree buffer on keep-alive power rail.
 *
 * Verilog wrapper for lpflow_clkbufkapwr with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkbufkapwr_4 (
    X    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkbufkapwr base (
        .X(X),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkbufkapwr: Clock tree buffer on keep-alive power rail.
 *
 * Verilog wrapper for lpflow_clkbufkapwr with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkbufkapwr_8 (
    X    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkbufkapwr base (
        .X(X),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkbufkapwr: Clock tree buffer on keep-alive power rail.
 *
 * Verilog wrapper for lpflow_clkbufkapwr with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkbufkapwr_16 (
    X    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkbufkapwr base (
        .X(X),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkinvkapwr: Clock tree inverter on keep-alive rail.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_clkinvkapwr: Clock tree inverter on keep-alive rail.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_clkinvkapwr (
    Y    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Y    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire not0_out_Y    ;
    wire pwrgood0_out_Y;

    //                                   Name      Output          Other arguments
    not                                  not0     (not0_out_Y    , A                      );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (pwrgood0_out_Y, not0_out_Y, KAPWR, VGND);
    buf                                  buf0     (Y             , pwrgood0_out_Y         );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_FUNCTIONAL_PP_V




































































 // FUNCTIONAL
























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkinvkapwr: Clock tree inverter on keep-alive rail.
 *
 * Verilog wrapper for lpflow_clkinvkapwr with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkinvkapwr_1 (
    Y    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Y    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkinvkapwr base (
        .Y(Y),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkinvkapwr: Clock tree inverter on keep-alive rail.
 *
 * Verilog wrapper for lpflow_clkinvkapwr with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkinvkapwr_2 (
    Y    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Y    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkinvkapwr base (
        .Y(Y),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkinvkapwr: Clock tree inverter on keep-alive rail.
 *
 * Verilog wrapper for lpflow_clkinvkapwr with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkinvkapwr_4 (
    Y    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Y    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkinvkapwr base (
        .Y(Y),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkinvkapwr: Clock tree inverter on keep-alive rail.
 *
 * Verilog wrapper for lpflow_clkinvkapwr with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkinvkapwr_8 (
    Y    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Y    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkinvkapwr base (
        .Y(Y),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_clkinvkapwr: Clock tree inverter on keep-alive rail.
 *
 * Verilog wrapper for lpflow_clkinvkapwr with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_clkinvkapwr_16 (
    Y    ,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Y    ;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_clkinvkapwr base (
        .Y(Y),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_decapkapwr: Decoupling capacitance filler on keep-alive
 *                    rail.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_decapkapwr: Decoupling capacitance filler on keep-alive
 *                    rail.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__lpflow_decapkapwr (
    VPWR ,
    KAPWR,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    input VPWR ;
    input KAPWR;
    input VGND ;
    input VPB  ;
    input VNB  ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_FUNCTIONAL_PP_V






















































 // FUNCTIONAL






























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_decapkapwr: Decoupling capacitance filler on keep-alive
 *                    rail.
 *
 * Verilog wrapper for lpflow_decapkapwr with size of 3 units
 * (invalid?).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_decapkapwr_3 (
    VPWR ,
    KAPWR,
    VGND ,
    VPB  ,
    VNB
);

    input VPWR ;
    input KAPWR;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__lpflow_decapkapwr base (
        .VPWR(VPWR),
        .KAPWR(KAPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/


















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_decapkapwr: Decoupling capacitance filler on keep-alive
 *                    rail.
 *
 * Verilog wrapper for lpflow_decapkapwr with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_decapkapwr_4 (
    VPWR ,
    KAPWR,
    VGND ,
    VPB  ,
    VNB
);

    input VPWR ;
    input KAPWR;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__lpflow_decapkapwr base (
        .VPWR(VPWR),
        .KAPWR(KAPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/


















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_decapkapwr: Decoupling capacitance filler on keep-alive
 *                    rail.
 *
 * Verilog wrapper for lpflow_decapkapwr with size of 6 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_decapkapwr_6 (
    VPWR ,
    KAPWR,
    VGND ,
    VPB  ,
    VNB
);

    input VPWR ;
    input KAPWR;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__lpflow_decapkapwr base (
        .VPWR(VPWR),
        .KAPWR(KAPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/


















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_decapkapwr: Decoupling capacitance filler on keep-alive
 *                    rail.
 *
 * Verilog wrapper for lpflow_decapkapwr with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_decapkapwr_8 (
    VPWR ,
    KAPWR,
    VGND ,
    VPB  ,
    VNB
);

    input VPWR ;
    input KAPWR;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__lpflow_decapkapwr base (
        .VPWR(VPWR),
        .KAPWR(KAPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/


















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_decapkapwr: Decoupling capacitance filler on keep-alive
 *                    rail.
 *
 * Verilog wrapper for lpflow_decapkapwr with size of 12 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_decapkapwr_12 (
    VPWR ,
    KAPWR,
    VGND ,
    VPB  ,
    VNB
);

    input VPWR ;
    input KAPWR;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hd__lpflow_decapkapwr base (
        .VPWR(VPWR),
        .KAPWR(KAPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/


















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputiso0n: Input isolator with inverted enable.
 *
 *                    X = (A & SLEEP_B)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_inputiso0n: Input isolator with inverted enable.
 *
 *                    X = (A & SLEEP_B)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_inputiso0n (
    X      ,
    A      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output X      ;
    input  A      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire and0_out_X;

    //                                   Name      Output      Other arguments
    and                                  and0     (and0_out_X, A, SLEEP_B            );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (X         , and0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_FUNCTIONAL_PP_V




































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputiso0n: Input isolator with inverted enable.
 *
 *                    X = (A & SLEEP_B)
 *
 * Verilog wrapper for lpflow_inputiso0n with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_inputiso0n_1 (
    X      ,
    A      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output X      ;
    input  A      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__lpflow_inputiso0n base (
        .X(X),
        .A(A),
        .SLEEP_B(SLEEP_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputiso0p: Input isolator with non-inverted enable.
 *
 *                    X = (A & !SLEEP_B)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_inputiso0p: Input isolator with non-inverted enable.
 *
 *                    X = (A & !SLEEP_B)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_inputiso0p (
    X    ,
    A    ,
    SLEEP,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  A    ;
    input  SLEEP;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire sleepn    ;
    wire and0_out_X;

    //                                   Name      Output      Other arguments
    not                                  not0     (sleepn    , SLEEP                 );
    and                                  and0     (and0_out_X, A, sleepn             );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (X         , and0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO0P_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO0P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputiso0p: Input isolator with non-inverted enable.
 *
 *                    X = (A & !SLEEP_B)
 *
 * Verilog wrapper for lpflow_inputiso0p with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_inputiso0p_1 (
    X    ,
    A    ,
    SLEEP,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  SLEEP;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_inputiso0p base (
        .X(X),
        .A(A),
        .SLEEP(SLEEP),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO0P_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputiso1n: Input isolation, inverted sleep.
 *
 *                    X = (A & SLEEP_B)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_inputiso1n: Input isolation, inverted sleep.
 *
 *                    X = (A & SLEEP_B)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_inputiso1n (
    X      ,
    A      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output X      ;
    input  A      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire SLEEP    ;
    wire or0_out_X;

    //                                   Name      Output     Other arguments
    not                                  not0     (SLEEP    , SLEEP_B              );
    or                                   or0      (or0_out_X, A, SLEEP             );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (X        , or0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputiso1n: Input isolation, inverted sleep.
 *
 *                    X = (A & SLEEP_B)
 *
 * Verilog wrapper for lpflow_inputiso1n with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_inputiso1n_1 (
    X      ,
    A      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output X      ;
    input  A      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__lpflow_inputiso1n base (
        .X(X),
        .A(A),
        .SLEEP_B(SLEEP_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputiso1p: Input isolation, noninverted sleep.
 *
 *                    X = (A & !SLEEP)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_inputiso1p: Input isolation, noninverted sleep.
 *
 *                    X = (A & !SLEEP)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_inputiso1p (
    X    ,
    A    ,
    SLEEP,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  A    ;
    input  SLEEP;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire or0_out_X;

    //                                   Name      Output     Other arguments
    or                                   or0      (or0_out_X, A, SLEEP             );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (X        , or0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_FUNCTIONAL_PP_V




































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputiso1p: Input isolation, noninverted sleep.
 *
 *                    X = (A & !SLEEP)
 *
 * Verilog wrapper for lpflow_inputiso1p with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_inputiso1p_1 (
    X    ,
    A    ,
    SLEEP,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  SLEEP;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_inputiso1p base (
        .X(X),
        .A(A),
        .SLEEP(SLEEP),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputisolatch: Latching input isolator with inverted enable.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_inputisolatch: Latching input isolator with inverted enable.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_inputisolatch (
    Q      ,
    D      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  D      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q;

    //                                     Name     Output  Other arguments
    sky130_fd_sc_hd__udp_dlatch$lP_pp$PG$N dlatch0 (buf_Q , D, SLEEP_B, 1'b0, VPWR, VGND);
    buf                                    buf0    (Q     , buf_Q                       );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_FUNCTIONAL_PP_V





































































 // FUNCTIONAL


































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_inputisolatch: Latching input isolator with inverted enable.
 *
 * Verilog wrapper for lpflow_inputisolatch with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_inputisolatch_1 (
    Q      ,
    D      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  D      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__lpflow_inputisolatch base (
        .Q(Q),
        .D(D),
        .SLEEP_B(SLEEP_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_isobufsrc: Input isolation, noninverted sleep.
 *
 *                   X = (!A | SLEEP)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_isobufsrc: Input isolation, noninverted sleep.
 *
 *                   X = (!A | SLEEP)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_isobufsrc (
    X    ,
    SLEEP,
    A    ,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  SLEEP;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire not0_out      ;
    wire and0_out_X    ;
    wire pwrgood0_out_X;

    //                                     Name      Output          Other arguments
    not                                    not0     (not0_out      , SLEEP                        );
    and                                    and0     (and0_out_X    , not0_out, A                  );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG$S pwrgood0 (pwrgood0_out_X, and0_out_X, VPWR, VGND, SLEEP);
    buf                                    buf0     (X             , pwrgood0_out_X               );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_isobufsrc: Input isolation, noninverted sleep.
 *
 *                   X = (!A | SLEEP)
 *
 * Verilog wrapper for lpflow_isobufsrc with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_isobufsrc_1 (
    X    ,
    SLEEP,
    A    ,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  SLEEP;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_isobufsrc base (
        .X(X),
        .SLEEP(SLEEP),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_isobufsrc: Input isolation, noninverted sleep.
 *
 *                   X = (!A | SLEEP)
 *
 * Verilog wrapper for lpflow_isobufsrc with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_isobufsrc_2 (
    X    ,
    SLEEP,
    A    ,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  SLEEP;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_isobufsrc base (
        .X(X),
        .SLEEP(SLEEP),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_isobufsrc: Input isolation, noninverted sleep.
 *
 *                   X = (!A | SLEEP)
 *
 * Verilog wrapper for lpflow_isobufsrc with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_isobufsrc_4 (
    X    ,
    SLEEP,
    A    ,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  SLEEP;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_isobufsrc base (
        .X(X),
        .SLEEP(SLEEP),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_isobufsrc: Input isolation, noninverted sleep.
 *
 *                   X = (!A | SLEEP)
 *
 * Verilog wrapper for lpflow_isobufsrc with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_isobufsrc_8 (
    X    ,
    SLEEP,
    A    ,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  SLEEP;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_isobufsrc base (
        .X(X),
        .SLEEP(SLEEP),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_isobufsrc: Input isolation, noninverted sleep.
 *
 *                   X = (!A | SLEEP)
 *
 * Verilog wrapper for lpflow_isobufsrc with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_isobufsrc_16 (
    X    ,
    SLEEP,
    A    ,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  SLEEP;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_isobufsrc base (
        .X(X),
        .SLEEP(SLEEP),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_isobufsrckapwr: Input isolation, noninverted sleep on
 *                        keep-alive power rail.
 *
 *                        X = (!A | SLEEP)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_isobufsrckapwr: Input isolation, noninverted sleep on
 *                        keep-alive power rail.
 *
 *                        X = (!A | SLEEP)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_isobufsrckapwr (
    X    ,
    SLEEP,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  SLEEP;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire not0_out       ;
    wire and0_out_X     ;
    wire pwrgood0_out_X ;
    wire pwrgood1_out_x2;

    //                                     Name      Output           Other arguments
    not                                    not0     (not0_out       , SLEEP                        );
    and                                    and0     (and0_out_X     , not0_out, A                  );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG$S pwrgood0 (pwrgood0_out_X , and0_out_X, VPWR, VGND, SLEEP);
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG   pwrgood1 (pwrgood1_out_x2, pwrgood0_out_X, KAPWR, VGND  );
    buf                                    buf0     (X              , pwrgood1_out_x2              );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_FUNCTIONAL_PP_V













































































 // FUNCTIONAL






































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_isobufsrckapwr: Input isolation, noninverted sleep on
 *                        keep-alive power rail.
 *
 *                        X = (!A | SLEEP)
 *
 * Verilog wrapper for lpflow_isobufsrckapwr with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 (
    X    ,
    SLEEP,
    A    ,
    KAPWR,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output X    ;
    input  SLEEP;
    input  A    ;
    input  KAPWR;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__lpflow_isobufsrckapwr base (
        .X(X),
        .SLEEP(SLEEP),
        .A(A),
        .KAPWR(KAPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_hl_isowell_tap: Level-shift buffer, low-to-high,
 *                                 isolated well on input buffer,
 *                                 vpb/vnb taps, double-row-height
 *                                 cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_lsbuf_lh_hl_isowell_tap: Level-shift buffer, low-to-high,
 *                                 isolated well on input buffer,
 *                                 vpb/vnb taps, double-row-height
 *                                 cell.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap (
    X     ,
    A     ,
    VPWRIN,
    VPWR  ,
    VGND  ,
    VPB
);

    // Module ports
    output X     ;
    input  A     ;
    input  VPWRIN;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;

    // Local signals
    wire pwrgood0_out_A;
    wire buf0_out_X    ;

    //                                   Name      Output          Other arguments
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (pwrgood0_out_A, A, VPWRIN, VGND       );
    buf                                  buf0     (buf0_out_X    , pwrgood0_out_A        );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood1 (X             , buf0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_FUNCTIONAL_PP_V





































































 // FUNCTIONAL




















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_hl_isowell_tap: Level-shift buffer, low-to-high,
 *                                 isolated well on input buffer,
 *                                 vpb/vnb taps, double-row-height
 *                                 cell.
 *
 * Verilog wrapper for lpflow_lsbuf_lh_hl_isowell_tap with
 * size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 (
    X     ,
    A     ,
    VPWRIN,
    VPWR  ,
    VGND  ,
    VPB
);

    output X     ;
    input  A     ;
    input  VPWRIN;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap base (
        .X(X),
        .A(A),
        .VPWRIN(VPWRIN),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_hl_isowell_tap: Level-shift buffer, low-to-high,
 *                                 isolated well on input buffer,
 *                                 vpb/vnb taps, double-row-height
 *                                 cell.
 *
 * Verilog wrapper for lpflow_lsbuf_lh_hl_isowell_tap with
 * size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 (
    X     ,
    A     ,
    VPWRIN,
    VPWR  ,
    VGND  ,
    VPB
);

    output X     ;
    input  A     ;
    input  VPWRIN;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap base (
        .X(X),
        .A(A),
        .VPWRIN(VPWRIN),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_hl_isowell_tap: Level-shift buffer, low-to-high,
 *                                 isolated well on input buffer,
 *                                 vpb/vnb taps, double-row-height
 *                                 cell.
 *
 * Verilog wrapper for lpflow_lsbuf_lh_hl_isowell_tap with
 * size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 (
    X     ,
    A     ,
    VPWRIN,
    VPWR  ,
    VGND  ,
    VPB
);

    output X     ;
    input  A     ;
    input  VPWRIN;
    input  VPWR  ;
    input  VGND  ;
    input  VPB   ;
    sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap base (
        .X(X),
        .A(A),
        .VPWRIN(VPWRIN),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_isowell: Level-shift buffer, low-to-high, isolated
 *                          well on input buffer, no taps,
 *                          double-row-height cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_lsbuf_lh_isowell: Level-shift buffer, low-to-high, isolated
 *                          well on input buffer, no taps,
 *                          double-row-height cell.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell (
    X       ,
    A       ,
    LOWLVPWR,
    VPWR    ,
    VGND    ,
    VPB     ,
    VNB
);

    // Module ports
    output X       ;
    input  A       ;
    input  LOWLVPWR;
    input  VPWR    ;
    input  VGND    ;
    input  VPB     ;
    input  VNB     ;

    // Local signals
    wire pwrgood0_out_A;
    wire buf0_out_X    ;

    //                                   Name      Output          Other arguments
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (pwrgood0_out_A, A, LOWLVPWR, VGND     );
    buf                                  buf0     (buf0_out_X    , pwrgood0_out_A        );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood1 (X             , buf0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_FUNCTIONAL_PP_V






































































 // FUNCTIONAL



















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_isowell: Level-shift buffer, low-to-high, isolated
 *                          well on input buffer, no taps,
 *                          double-row-height cell.
 *
 * Verilog wrapper for lpflow_lsbuf_lh_isowell with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 (
    X       ,
    A       ,
    LOWLVPWR,
    VPWR    ,
    VGND    ,
    VPB     ,
    VNB
);

    output X       ;
    input  A       ;
    input  LOWLVPWR;
    input  VPWR    ;
    input  VGND    ;
    input  VPB     ;
    input  VNB     ;
    sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell base (
        .X(X),
        .A(A),
        .LOWLVPWR(LOWLVPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_isowell_tap: Level-shift buffer, low-to-high,
 *                              isolated well on input buffer, vpb/vnb
 *                              taps, double-row-height cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lpflow_lsbuf_lh_isowell_tap: Level-shift buffer, low-to-high,
 *                              isolated well on input buffer, vpb/vnb
 *                              taps, double-row-height cell.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap (
    X       ,
    A       ,
    LOWLVPWR,
    VPWR    ,
    VGND    ,
    VPB
);

    // Module ports
    output X       ;
    input  A       ;
    input  LOWLVPWR;
    input  VPWR    ;
    input  VGND    ;
    input  VPB     ;

    // Local signals
    wire pwrgood0_out_A;
    wire buf0_out_X    ;

    //                                   Name      Output          Other arguments
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood0 (pwrgood0_out_A, A, LOWLVPWR, VGND     );
    buf                                  buf0     (buf0_out_X    , pwrgood0_out_A        );
    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG pwrgood1 (X             , buf0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_FUNCTIONAL_PP_V




































































 // FUNCTIONAL


















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_isowell_tap: Level-shift buffer, low-to-high,
 *                              isolated well on input buffer, vpb/vnb
 *                              taps, double-row-height cell.
 *
 * Verilog wrapper for lpflow_lsbuf_lh_isowell_tap with
 * size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 (
    X       ,
    A       ,
    LOWLVPWR,
    VPWR    ,
    VGND    ,
    VPB
);

    output X       ;
    input  A       ;
    input  LOWLVPWR;
    input  VPWR    ;
    input  VGND    ;
    input  VPB     ;
    sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap base (
        .X(X),
        .A(A),
        .LOWLVPWR(LOWLVPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_isowell_tap: Level-shift buffer, low-to-high,
 *                              isolated well on input buffer, vpb/vnb
 *                              taps, double-row-height cell.
 *
 * Verilog wrapper for lpflow_lsbuf_lh_isowell_tap with
 * size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 (
    X       ,
    A       ,
    LOWLVPWR,
    VPWR    ,
    VGND    ,
    VPB
);

    output X       ;
    input  A       ;
    input  LOWLVPWR;
    input  VPWR    ;
    input  VGND    ;
    input  VPB     ;
    sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap base (
        .X(X),
        .A(A),
        .LOWLVPWR(LOWLVPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lpflow_lsbuf_lh_isowell_tap: Level-shift buffer, low-to-high,
 *                              isolated well on input buffer, vpb/vnb
 *                              taps, double-row-height cell.
 *
 * Verilog wrapper for lpflow_lsbuf_lh_isowell_tap with
 * size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 (
    X       ,
    A       ,
    LOWLVPWR,
    VPWR    ,
    VGND    ,
    VPB
);

    output X       ;
    input  A       ;
    input  LOWLVPWR;
    input  VPWR    ;
    input  VGND    ;
    input  VPB     ;
    sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap base (
        .X(X),
        .A(A),
        .LOWLVPWR(LOWLVPWR),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * macro_sparecell: Macro cell for metal-mask-only revisioning,
 *                  containing inverter, 2-input NOR, 2-input NAND,
 *                  and constant cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * macro_sparecell: Macro cell for metal-mask-only revisioning,
 *                  containing inverter, 2-input NOR, 2-input NAND,
 *                  and constant cell.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import sub cells.

`celldefine
module sky130_fd_sc_hd__macro_sparecell (
    LO  ,
    VGND,
    VNB ,
    VPB ,
    VPWR
);

    // Module ports
    output LO  ;
    input  VGND;
    input  VNB ;
    input  VPB ;
    input  VPWR;

    // Local signals
    wire nor2left ;
    wire invleft  ;
    wire nor2right;
    wire invright ;
    wire nd2left  ;
    wire nd2right ;
    wire tielo    ;
    wire net7     ;

    //                       Name    Output         Other arguments
    sky130_fd_sc_hd__inv_2   inv0   (.A(nor2left) , .Y(invleft), .VPWR(VPWR), .VGND(VGND), .VNB(VNB), .VPB(VPB)                );
    sky130_fd_sc_hd__inv_2   inv1   (.A(nor2right), .Y(invright), .VPWR(VPWR), .VGND(VGND), .VNB(VNB), .VPB(VPB)               );
    sky130_fd_sc_hd__nor2_2  nor20  (.B(nd2left)  , .A(nd2left), .Y(nor2left), .VPWR(VPWR), .VGND(VGND), .VNB(VNB), .VPB(VPB)  );
    sky130_fd_sc_hd__nor2_2  nor21  (.B(nd2right) , .A(nd2right), .Y(nor2right), .VPWR(VPWR), .VGND(VGND), .VNB(VNB), .VPB(VPB));
    sky130_fd_sc_hd__nand2_2 nand20 (.B(tielo)    , .A(tielo), .Y(nd2right), .VPWR(VPWR), .VGND(VGND), .VNB(VNB), .VPB(VPB)    );
    sky130_fd_sc_hd__nand2_2 nand21 (.B(tielo)    , .A(tielo), .Y(nd2left), .VPWR(VPWR), .VGND(VGND), .VNB(VNB), .VPB(VPB)     );
    sky130_fd_sc_hd__conb_1  conb0  (.LO(tielo)   , .HI(net7), .VPWR(VPWR), .VGND(VGND), .VNB(VNB), .VPB(VPB)                  );
    buf                      buf0   (LO           , tielo                                                                      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__MACRO_SPARECELL_FUNCTIONAL_PP_V













































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MACRO_SPARECELL_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * maj3: 3-input majority vote.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * maj3: 3-input majority vote.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__maj3 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire and0_out         ;
    wire and1_out         ;
    wire or1_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , B, A                 );
    and                                and0        (and0_out         , or0_out, C           );
    and                                and1        (and1_out         , A, B                 );
    or                                 or1         (or1_out_X        , and1_out, and0_out   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or1_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__MAJ3_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MAJ3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * maj3: 3-input majority vote.
 *
 * Verilog wrapper for maj3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__maj3_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__maj3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MAJ3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * maj3: 3-input majority vote.
 *
 * Verilog wrapper for maj3 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__maj3_2 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__maj3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MAJ3_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * maj3: 3-input majority vote.
 *
 * Verilog wrapper for maj3 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__maj3_4 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__maj3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MAJ3_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2: 2-input multiplexer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * mux2: 2-input multiplexer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__mux2 (
    X   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire mux_2to10_out_X  ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    sky130_fd_sc_hd__udp_mux_2to1      mux_2to10   (mux_2to10_out_X  , A0, A1, S                  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, mux_2to10_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2_FUNCTIONAL_PP_V






































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2: 2-input multiplexer.
 *
 * Verilog wrapper for mux2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux2_1 (
    X   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux2 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .S(S),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2: 2-input multiplexer.
 *
 * Verilog wrapper for mux2 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux2_2 (
    X   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux2 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .S(S),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2: 2-input multiplexer.
 *
 * Verilog wrapper for mux2 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux2_4 (
    X   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux2 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .S(S),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2: 2-input multiplexer.
 *
 * Verilog wrapper for mux2 with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux2_8 (
    X   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux2 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .S(S),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2i: 2-input multiplexer, output inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * mux2i: 2-input multiplexer, output inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__mux2i (
    Y   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire mux_2to1_n0_out_Y;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    sky130_fd_sc_hd__udp_mux_2to1_N    mux_2to1_n0 (mux_2to1_n0_out_Y, A0, A1, S                    );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, mux_2to1_n0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y            );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2I_FUNCTIONAL_PP_V






































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2I_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2i: 2-input multiplexer, output inverted.
 *
 * Verilog wrapper for mux2i with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux2i_1 (
    Y   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux2i base (
        .Y(Y),
        .A0(A0),
        .A1(A1),
        .S(S),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2I_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2i: 2-input multiplexer, output inverted.
 *
 * Verilog wrapper for mux2i with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux2i_2 (
    Y   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux2i base (
        .Y(Y),
        .A0(A0),
        .A1(A1),
        .S(S),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2I_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2i: 2-input multiplexer, output inverted.
 *
 * Verilog wrapper for mux2i with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux2i_4 (
    Y   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux2i base (
        .Y(Y),
        .A0(A0),
        .A1(A1),
        .S(S),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX2I_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux4: 4-input multiplexer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * mux4: 4-input multiplexer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__mux4 (
    X   ,
    A0  ,
    A1  ,
    A2  ,
    A3  ,
    S0  ,
    S1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A0  ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  S0  ;
    input  S1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire mux_4to20_out_X  ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    sky130_fd_sc_hd__udp_mux_4to2      mux_4to20   (mux_4to20_out_X  , A0, A1, A2, A3, S0, S1     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, mux_4to20_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__MUX4_FUNCTIONAL_PP_V












































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux4: 4-input multiplexer.
 *
 * Verilog wrapper for mux4 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux4_1 (
    X   ,
    A0  ,
    A1  ,
    A2  ,
    A3  ,
    S0  ,
    S1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  S0  ;
    input  S1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux4 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .S0(S0),
        .S1(S1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX4_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux4: 4-input multiplexer.
 *
 * Verilog wrapper for mux4 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux4_2 (
    X   ,
    A0  ,
    A1  ,
    A2  ,
    A3  ,
    S0  ,
    S1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  S0  ;
    input  S1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux4 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .S0(S0),
        .S1(S1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX4_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux4: 4-input multiplexer.
 *
 * Verilog wrapper for mux4 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__mux4_4 (
    X   ,
    A0  ,
    A1  ,
    A2  ,
    A3  ,
    S0  ,
    S1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  S0  ;
    input  S1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__mux4 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .S0(S0),
        .S1(S1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__MUX4_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2: 2-input NAND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand2: 2-input NAND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nand2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out_Y      , B, A                   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2: 2-input NAND.
 *
 * Verilog wrapper for nand2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand2_1 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2: 2-input NAND.
 *
 * Verilog wrapper for nand2 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand2_2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2: 2-input NAND.
 *
 * Verilog wrapper for nand2 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand2_4 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2: 2-input NAND.
 *
 * Verilog wrapper for nand2 with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand2_8 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2b: 2-input NAND, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand2b: 2-input NAND, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nand2b (
    Y   ,
    A_N ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A_N ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire or0_out_Y        ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , B                    );
    or                                 or0         (or0_out_Y        , not0_out, A_N        );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, or0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2B_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2b: 2-input NAND, first input inverted.
 *
 * Verilog wrapper for nand2b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand2b_1 (
    Y   ,
    A_N ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand2b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2b: 2-input NAND, first input inverted.
 *
 * Verilog wrapper for nand2b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand2b_2 (
    Y   ,
    A_N ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand2b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2b: 2-input NAND, first input inverted.
 *
 * Verilog wrapper for nand2b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand2b_4 (
    Y   ,
    A_N ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand2b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND2B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3: 3-input NAND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand3: 3-input NAND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nand3 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out_Y      , B, A, C                );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3: 3-input NAND.
 *
 * Verilog wrapper for nand3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand3_1 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand3 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3: 3-input NAND.
 *
 * Verilog wrapper for nand3 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand3_2 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand3 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3: 3-input NAND.
 *
 * Verilog wrapper for nand3 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand3_4 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand3 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3b: 3-input NAND, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand3b: 3-input NAND, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nand3b (
    Y   ,
    A_N ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , A_N                    );
    nand                               nand0       (nand0_out_Y      , B, not0_out, C         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3B_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3b: 3-input NAND, first input inverted.
 *
 * Verilog wrapper for nand3b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand3b_1 (
    Y   ,
    A_N ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand3b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3b: 3-input NAND, first input inverted.
 *
 * Verilog wrapper for nand3b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand3b_2 (
    Y   ,
    A_N ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand3b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3b: 3-input NAND, first input inverted.
 *
 * Verilog wrapper for nand3b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand3b_4 (
    Y   ,
    A_N ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand3b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND3B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4: 4-input NAND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand4: 4-input NAND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nand4 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out_Y      , D, C, B, A             );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4: 4-input NAND.
 *
 * Verilog wrapper for nand4 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4_1 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4: 4-input NAND.
 *
 * Verilog wrapper for nand4 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4_2 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4: 4-input NAND.
 *
 * Verilog wrapper for nand4 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4_4 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4b: 4-input NAND, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand4b: 4-input NAND, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nand4b (
    Y   ,
    A_N ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , A_N                    );
    nand                               nand0       (nand0_out_Y      , D, C, B, not0_out      );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4B_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4b: 4-input NAND, first input inverted.
 *
 * Verilog wrapper for nand4b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4b_1 (
    Y   ,
    A_N ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4b: 4-input NAND, first input inverted.
 *
 * Verilog wrapper for nand4b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4b_2 (
    Y   ,
    A_N ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4b: 4-input NAND, first input inverted.
 *
 * Verilog wrapper for nand4b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4b_4 (
    Y   ,
    A_N ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4b base (
        .Y(Y),
        .A_N(A_N),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4bb: 4-input NAND, first two inputs inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand4bb: 4-input NAND, first two inputs inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nand4bb (
    Y   ,
    A_N ,
    B_N ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A_N ;
    input  B_N ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire or0_out_Y        ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out        , D, C                 );
    or                                 or0         (or0_out_Y        , B_N, A_N, nand0_out  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, or0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4BB_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4BB_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4bb: 4-input NAND, first two inputs inverted.
 *
 * Verilog wrapper for nand4bb with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4bb_1 (
    Y   ,
    A_N ,
    B_N ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B_N ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4bb base (
        .Y(Y),
        .A_N(A_N),
        .B_N(B_N),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4BB_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4bb: 4-input NAND, first two inputs inverted.
 *
 * Verilog wrapper for nand4bb with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4bb_2 (
    Y   ,
    A_N ,
    B_N ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B_N ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4bb base (
        .Y(Y),
        .A_N(A_N),
        .B_N(B_N),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4BB_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand4bb: 4-input NAND, first two inputs inverted.
 *
 * Verilog wrapper for nand4bb with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nand4bb_4 (
    Y   ,
    A_N ,
    B_N ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A_N ;
    input  B_N ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nand4bb base (
        .Y(Y),
        .A_N(A_N),
        .B_N(B_N),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NAND4BB_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2: 2-input NOR.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor2: 2-input NOR.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nor2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out_Y       , A, B                  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2: 2-input NOR.
 *
 * Verilog wrapper for nor2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor2_1 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2: 2-input NOR.
 *
 * Verilog wrapper for nor2 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor2_2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2: 2-input NOR.
 *
 * Verilog wrapper for nor2 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor2_4 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2: 2-input NOR.
 *
 * Verilog wrapper for nor2 with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor2_8 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2b: 2-input NOR, first input inverted.
 *
 *        Y = !(A | B | C | !D)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor2b: 2-input NOR, first input inverted.
 *
 *        Y = !(A | B | C | !D)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nor2b (
    Y   ,
    A   ,
    B_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire and0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , A                     );
    and                                and0        (and0_out_Y       , not0_out, B_N         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, and0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2B_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2b: 2-input NOR, first input inverted.
 *
 *        Y = !(A | B | C | !D)
 *
 * Verilog wrapper for nor2b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor2b_1 (
    Y   ,
    A   ,
    B_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor2b base (
        .Y(Y),
        .A(A),
        .B_N(B_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2b: 2-input NOR, first input inverted.
 *
 *        Y = !(A | B | C | !D)
 *
 * Verilog wrapper for nor2b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor2b_2 (
    Y   ,
    A   ,
    B_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor2b base (
        .Y(Y),
        .A(A),
        .B_N(B_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2b: 2-input NOR, first input inverted.
 *
 *        Y = !(A | B | C | !D)
 *
 * Verilog wrapper for nor2b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor2b_4 (
    Y   ,
    A   ,
    B_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor2b base (
        .Y(Y),
        .A(A),
        .B_N(B_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR2B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3: 3-input NOR.
 *
 *       Y = !(A | B | C | !D)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor3: 3-input NOR.
 *
 *       Y = !(A | B | C | !D)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nor3 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out_Y       , C, A, B               );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3: 3-input NOR.
 *
 *       Y = !(A | B | C | !D)
 *
 * Verilog wrapper for nor3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor3_1 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor3 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3: 3-input NOR.
 *
 *       Y = !(A | B | C | !D)
 *
 * Verilog wrapper for nor3 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor3_2 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor3 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3: 3-input NOR.
 *
 *       Y = !(A | B | C | !D)
 *
 * Verilog wrapper for nor3 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor3_4 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor3 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3b: 3-input NOR, first input inverted.
 *
 *        Y = (!(A | B)) & !C)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor3b: 3-input NOR, first input inverted.
 *
 *        Y = (!(A | B)) & !C)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nor3b (
    Y   ,
    A   ,
    B   ,
    C_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out         ;
    wire and0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out         , A, B                  );
    and                                and0        (and0_out_Y       , C_N, nor0_out         );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, and0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3B_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3b: 3-input NOR, first input inverted.
 *
 *        Y = (!(A | B)) & !C)
 *
 * Verilog wrapper for nor3b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor3b_1 (
    Y   ,
    A   ,
    B   ,
    C_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor3b base (
        .Y(Y),
        .A(A),
        .B(B),
        .C_N(C_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3b: 3-input NOR, first input inverted.
 *
 *        Y = (!(A | B)) & !C)
 *
 * Verilog wrapper for nor3b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor3b_2 (
    Y   ,
    A   ,
    B   ,
    C_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor3b base (
        .Y(Y),
        .A(A),
        .B(B),
        .C_N(C_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3b: 3-input NOR, first input inverted.
 *
 *        Y = (!(A | B)) & !C)
 *
 * Verilog wrapper for nor3b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor3b_4 (
    Y   ,
    A   ,
    B   ,
    C_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor3b base (
        .Y(Y),
        .A(A),
        .B(B),
        .C_N(C_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR3B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4: 4-input NOR.
 *
 *       Y = !(A | B | C | D)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor4: 4-input NOR.
 *
 *       Y = !(A | B | C | D)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nor4 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out_Y       , A, B, C, D            );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4: 4-input NOR.
 *
 *       Y = !(A | B | C | D)
 *
 * Verilog wrapper for nor4 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4_1 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4: 4-input NOR.
 *
 *       Y = !(A | B | C | D)
 *
 * Verilog wrapper for nor4 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4_2 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4: 4-input NOR.
 *
 *       Y = !(A | B | C | D)
 *
 * Verilog wrapper for nor4 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4_4 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4b: 4-input NOR, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor4b: 4-input NOR, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nor4b (
    Y   ,
    A   ,
    B   ,
    C   ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , D_N                   );
    nor                                nor0        (nor0_out_Y       , A, B, C, not0_out     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4B_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4b: 4-input NOR, first input inverted.
 *
 * Verilog wrapper for nor4b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4b_1 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4b base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4b: 4-input NOR, first input inverted.
 *
 * Verilog wrapper for nor4b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4b_2 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4b base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4b: 4-input NOR, first input inverted.
 *
 * Verilog wrapper for nor4b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4b_4 (
    Y   ,
    A   ,
    B   ,
    C   ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4b base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4bb: 4-input NOR, first two inputs inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor4bb: 4-input NOR, first two inputs inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__nor4bb (
    Y   ,
    A   ,
    B   ,
    C_N ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out         ;
    wire and0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out         , A, B                  );
    and                                and0        (and0_out_Y       , nor0_out, C_N, D_N    );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, and0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4BB_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4BB_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4bb: 4-input NOR, first two inputs inverted.
 *
 * Verilog wrapper for nor4bb with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4bb_1 (
    Y   ,
    A   ,
    B   ,
    C_N ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4bb base (
        .Y(Y),
        .A(A),
        .B(B),
        .C_N(C_N),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4BB_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4bb: 4-input NOR, first two inputs inverted.
 *
 * Verilog wrapper for nor4bb with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4bb_2 (
    Y   ,
    A   ,
    B   ,
    C_N ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4bb base (
        .Y(Y),
        .A(A),
        .B(B),
        .C_N(C_N),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4BB_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor4bb: 4-input NOR, first two inputs inverted.
 *
 * Verilog wrapper for nor4bb with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__nor4bb_4 (
    Y   ,
    A   ,
    B   ,
    C_N ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__nor4bb base (
        .Y(Y),
        .A(A),
        .B(B),
        .C_N(C_N),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__NOR4BB_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2bb2a: 2-input NAND and 2-input OR into 2-input AND.
 *
 *         X = (!(A1 & A2) & (B1 | B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o2bb2a: 2-input NAND and 2-input OR into 2-input AND.
 *
 *         X = (!(A1 & A2) & (B1 | B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o2bb2a (
    X   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire or0_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out        , A2_N, A1_N            );
    or                                 or0         (or0_out          , B2, B1                );
    and                                and0        (and0_out_X       , nand0_out, or0_out    );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2A_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2bb2a: 2-input NAND and 2-input OR into 2-input AND.
 *
 *         X = (!(A1 & A2) & (B1 | B2))
 *
 * Verilog wrapper for o2bb2a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2bb2a_1 (
    X   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2bb2a base (
        .X(X),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2bb2a: 2-input NAND and 2-input OR into 2-input AND.
 *
 *         X = (!(A1 & A2) & (B1 | B2))
 *
 * Verilog wrapper for o2bb2a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2bb2a_2 (
    X   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2bb2a base (
        .X(X),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2bb2a: 2-input NAND and 2-input OR into 2-input AND.
 *
 *         X = (!(A1 & A2) & (B1 | B2))
 *
 * Verilog wrapper for o2bb2a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2bb2a_4 (
    X   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2bb2a base (
        .X(X),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2bb2ai: 2-input NAND and 2-input OR into 2-input NAND.
 *
 *          Y = !(!(A1 & A2) & (B1 | B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o2bb2ai: 2-input NAND and 2-input OR into 2-input NAND.
 *
 *          Y = !(!(A1 & A2) & (B1 | B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o2bb2ai (
    Y   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire or0_out          ;
    wire nand1_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out        , A2_N, A1_N             );
    or                                 or0         (or0_out          , B2, B1                 );
    nand                               nand1       (nand1_out_Y      , nand0_out, or0_out     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand1_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2AI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2bb2ai: 2-input NAND and 2-input OR into 2-input NAND.
 *
 *          Y = !(!(A1 & A2) & (B1 | B2))
 *
 * Verilog wrapper for o2bb2ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2bb2ai_1 (
    Y   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2bb2ai base (
        .Y(Y),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2bb2ai: 2-input NAND and 2-input OR into 2-input NAND.
 *
 *          Y = !(!(A1 & A2) & (B1 | B2))
 *
 * Verilog wrapper for o2bb2ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2bb2ai_2 (
    Y   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2bb2ai base (
        .Y(Y),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2bb2ai: 2-input NAND and 2-input OR into 2-input NAND.
 *
 *          Y = !(!(A1 & A2) & (B1 | B2))
 *
 * Verilog wrapper for o2bb2ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2bb2ai_4 (
    Y   ,
    A1_N,
    A2_N,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1_N;
    input  A2_N;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2bb2ai base (
        .Y(Y),
        .A1_N(A1_N),
        .A2_N(A2_N),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2BB2AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21a: 2-input OR into first input of 2-input AND.
 *
 *       X = ((A1 | A2) & B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o21a: 2-input OR into first input of 2-input AND.
 *
 *       X = ((A1 | A2) & B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o21a (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1                );
    and                                and0        (and0_out_X       , or0_out, B1           );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O21A_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21a: 2-input OR into first input of 2-input AND.
 *
 *       X = ((A1 | A2) & B1)
 *
 * Verilog wrapper for o21a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21a_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21a: 2-input OR into first input of 2-input AND.
 *
 *       X = ((A1 | A2) & B1)
 *
 * Verilog wrapper for o21a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21a_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21a: 2-input OR into first input of 2-input AND.
 *
 *       X = ((A1 | A2) & B1)
 *
 * Verilog wrapper for o21a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21a_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o21ai (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1                 );
    nand                               nand0       (nand0_out_Y      , B1, or0_out            );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O21AI_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog wrapper for o21ai with size of 0 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21ai_0 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21AI_0_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog wrapper for o21ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21ai_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog wrapper for o21ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21ai_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog wrapper for o21ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21ai_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ba: 2-input OR into first input of 2-input AND,
 *        2nd input inverted.
 *
 *        X = ((A1 | A2) & !B1_N)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o21ba: 2-input OR into first input of 2-input AND,
 *        2nd input inverted.
 *
 *        X = ((A1 | A2) & !B1_N)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o21ba (
    X   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out         ;
    wire nor1_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out         , A1, A2                );
    nor                                nor1        (nor1_out_X       , B1_N, nor0_out        );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, nor1_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O21BA_FUNCTIONAL_PP_V











































































 // FUNCTIONAL









































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21BA_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ba: 2-input OR into first input of 2-input AND,
 *        2nd input inverted.
 *
 *        X = ((A1 | A2) & !B1_N)
 *
 * Verilog wrapper for o21ba with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21ba_1 (
    X   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21ba base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21BA_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ba: 2-input OR into first input of 2-input AND,
 *        2nd input inverted.
 *
 *        X = ((A1 | A2) & !B1_N)
 *
 * Verilog wrapper for o21ba with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21ba_2 (
    X   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21ba base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21BA_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ba: 2-input OR into first input of 2-input AND,
 *        2nd input inverted.
 *
 *        X = ((A1 | A2) & !B1_N)
 *
 * Verilog wrapper for o21ba with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21ba_4 (
    X   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21ba base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21BA_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21bai: 2-input OR into first input of 2-input NAND, 2nd iput
 *         inverted.
 *
 *         Y = !((A1 | A2) & !B1_N)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o21bai: 2-input OR into first input of 2-input NAND, 2nd iput
 *         inverted.
 *
 *         Y = !((A1 | A2) & !B1_N)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o21bai (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire b                ;
    wire or0_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    not                                not0        (b                , B1_N                   );
    or                                 or0         (or0_out          , A2, A1                 );
    nand                               nand0       (nand0_out_Y      , b, or0_out             );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O21BAI_FUNCTIONAL_PP_V













































































 // FUNCTIONAL













































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21BAI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21bai: 2-input OR into first input of 2-input NAND, 2nd iput
 *         inverted.
 *
 *         Y = !((A1 | A2) & !B1_N)
 *
 * Verilog wrapper for o21bai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21bai_1 (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21bai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21BAI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21bai: 2-input OR into first input of 2-input NAND, 2nd iput
 *         inverted.
 *
 *         Y = !((A1 | A2) & !B1_N)
 *
 * Verilog wrapper for o21bai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21bai_2 (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21bai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21BAI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21bai: 2-input OR into first input of 2-input NAND, 2nd iput
 *         inverted.
 *
 *         Y = !((A1 | A2) & !B1_N)
 *
 * Verilog wrapper for o21bai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o21bai_4 (
    Y   ,
    A1  ,
    A2  ,
    B1_N,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1_N;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o21bai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1_N(B1_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O21BAI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22a: 2-input OR into both inputs of 2-input AND.
 *
 *       X = ((A1 | A2) & (B1 | B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o22a: 2-input OR into both inputs of 2-input AND.
 *
 *       X = ((A1 | A2) & (B1 | B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o22a (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire or1_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1                );
    or                                 or1         (or1_out          , B2, B1                );
    and                                and0        (and0_out_X       , or0_out, or1_out      );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O22A_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O22A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22a: 2-input OR into both inputs of 2-input AND.
 *
 *       X = ((A1 | A2) & (B1 | B2))
 *
 * Verilog wrapper for o22a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o22a_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o22a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O22A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22a: 2-input OR into both inputs of 2-input AND.
 *
 *       X = ((A1 | A2) & (B1 | B2))
 *
 * Verilog wrapper for o22a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o22a_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o22a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O22A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22a: 2-input OR into both inputs of 2-input AND.
 *
 *       X = ((A1 | A2) & (B1 | B2))
 *
 * Verilog wrapper for o22a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o22a_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o22a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O22A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22ai: 2-input OR into both inputs of 2-input NAND.
 *
 *        Y = !((A1 | A2) & (B1 | B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o22ai: 2-input OR into both inputs of 2-input NAND.
 *
 *        Y = !((A1 | A2) & (B1 | B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o22ai (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out         ;
    wire nor1_out         ;
    wire or0_out_Y        ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out         , B1, B2               );
    nor                                nor1        (nor1_out         , A1, A2               );
    or                                 or0         (or0_out_Y        , nor1_out, nor0_out   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, or0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O22AI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O22AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22ai: 2-input OR into both inputs of 2-input NAND.
 *
 *        Y = !((A1 | A2) & (B1 | B2))
 *
 * Verilog wrapper for o22ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o22ai_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o22ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O22AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22ai: 2-input OR into both inputs of 2-input NAND.
 *
 *        Y = !((A1 | A2) & (B1 | B2))
 *
 * Verilog wrapper for o22ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o22ai_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o22ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O22AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22ai: 2-input OR into both inputs of 2-input NAND.
 *
 *        Y = !((A1 | A2) & (B1 | B2))
 *
 * Verilog wrapper for o22ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o22ai_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o22ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O22AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o31a: 3-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o31a: 3-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o31a (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1, A3            );
    and                                and0        (and0_out_X       , or0_out, B1           );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O31A_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O31A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o31a: 3-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & B1)
 *
 * Verilog wrapper for o31a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o31a_1 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o31a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O31A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o31a: 3-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & B1)
 *
 * Verilog wrapper for o31a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o31a_2 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o31a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O31A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o31a: 3-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & B1)
 *
 * Verilog wrapper for o31a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o31a_4 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o31a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O31A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o31ai: 3-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o31ai: 3-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o31ai (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1, A3             );
    nand                               nand0       (nand0_out_Y      , B1, or0_out            );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O31AI_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O31AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o31ai: 3-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & B1)
 *
 * Verilog wrapper for o31ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o31ai_1 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o31ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O31AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o31ai: 3-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & B1)
 *
 * Verilog wrapper for o31ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o31ai_2 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o31ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O31AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o31ai: 3-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & B1)
 *
 * Verilog wrapper for o31ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o31ai_4 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o31ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O31AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o32a: 3-input OR and 2-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o32a: 3-input OR and 2-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o32a (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire or1_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1, A3            );
    or                                 or1         (or1_out          , B2, B1                );
    and                                and0        (and0_out_X       , or0_out, or1_out      );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O32A_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL



















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O32A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o32a: 3-input OR and 2-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog wrapper for o32a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o32a_1 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o32a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O32A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o32a: 3-input OR and 2-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog wrapper for o32a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o32a_2 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o32a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O32A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o32a: 3-input OR and 2-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog wrapper for o32a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o32a_4 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o32a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O32A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o32ai: 3-input OR and 2-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o32ai: 3-input OR and 2-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o32ai (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out         ;
    wire nor1_out         ;
    wire or0_out_Y        ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    nor                                nor0        (nor0_out         , A3, A1, A2           );
    nor                                nor1        (nor1_out         , B1, B2               );
    or                                 or0         (or0_out_Y        , nor1_out, nor0_out   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, or0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O32AI_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL



















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O32AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o32ai: 3-input OR and 2-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog wrapper for o32ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o32ai_1 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o32ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O32AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o32ai: 3-input OR and 2-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog wrapper for o32ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o32ai_2 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o32ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O32AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o32ai: 3-input OR and 2-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3) & (B1 | B2))
 *
 * Verilog wrapper for o32ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o32ai_4 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o32ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O32AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o41a: 4-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o41a: 4-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o41a (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A4, A3, A2, A1        );
    and                                and0        (and0_out_X       , or0_out, B1           );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O41A_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O41A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o41a: 4-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog wrapper for o41a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o41a_1 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o41a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O41A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o41a: 4-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog wrapper for o41a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o41a_2 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o41a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O41A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o41a: 4-input OR into 2-input AND.
 *
 *       X = ((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog wrapper for o41a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o41a_4 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o41a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O41A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o41ai: 4-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o41ai: 4-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o41ai (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A4, A3, A2, A1         );
    nand                               nand0       (nand0_out_Y      , B1, or0_out            );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O41AI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O41AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o41ai: 4-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog wrapper for o41ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o41ai_1 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o41ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O41AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o41ai: 4-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog wrapper for o41ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o41ai_2 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o41ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O41AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o41ai: 4-input OR into 2-input NAND.
 *
 *        Y = !((A1 | A2 | A3 | A4) & B1)
 *
 * Verilog wrapper for o41ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o41ai_4 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    A4  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  A4  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o41ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .A4(A4),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O41AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o211a: 2-input OR into first input of 3-input AND.
 *
 *        X = ((A1 | A2) & B1 & C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o211a: 2-input OR into first input of 3-input AND.
 *
 *        X = ((A1 | A2) & B1 & C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o211a (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1                );
    and                                and0        (and0_out_X       , or0_out, B1, C1       );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O211A_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O211A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o211a: 2-input OR into first input of 3-input AND.
 *
 *        X = ((A1 | A2) & B1 & C1)
 *
 * Verilog wrapper for o211a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o211a_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o211a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O211A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o211a: 2-input OR into first input of 3-input AND.
 *
 *        X = ((A1 | A2) & B1 & C1)
 *
 * Verilog wrapper for o211a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o211a_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o211a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O211A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o211a: 2-input OR into first input of 3-input AND.
 *
 *        X = ((A1 | A2) & B1 & C1)
 *
 * Verilog wrapper for o211a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o211a_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o211a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O211A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o211ai: 2-input OR into first input of 3-input NAND.
 *
 *         Y = !((A1 | A2) & B1 & C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o211ai: 2-input OR into first input of 3-input NAND.
 *
 *         Y = !((A1 | A2) & B1 & C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o211ai (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1                 );
    nand                               nand0       (nand0_out_Y      , C1, or0_out, B1        );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O211AI_FUNCTIONAL_PP_V












































































 // FUNCTIONAL











































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O211AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o211ai: 2-input OR into first input of 3-input NAND.
 *
 *         Y = !((A1 | A2) & B1 & C1)
 *
 * Verilog wrapper for o211ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o211ai_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o211ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O211AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o211ai: 2-input OR into first input of 3-input NAND.
 *
 *         Y = !((A1 | A2) & B1 & C1)
 *
 * Verilog wrapper for o211ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o211ai_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o211ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O211AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o211ai: 2-input OR into first input of 3-input NAND.
 *
 *         Y = !((A1 | A2) & B1 & C1)
 *
 * Verilog wrapper for o211ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o211ai_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o211ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O211AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o221a: 2-input OR into first two inputs of 3-input AND.
 *
 *        X = ((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o221a: 2-input OR into first two inputs of 3-input AND.
 *
 *        X = ((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o221a (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire or1_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , B2, B1                );
    or                                 or1         (or1_out          , A2, A1                );
    and                                and0        (and0_out_X       , or0_out, or1_out, C1  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O221A_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL



















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O221A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o221a: 2-input OR into first two inputs of 3-input AND.
 *
 *        X = ((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog wrapper for o221a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o221a_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o221a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O221A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o221a: 2-input OR into first two inputs of 3-input AND.
 *
 *        X = ((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog wrapper for o221a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o221a_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o221a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O221A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o221a: 2-input OR into first two inputs of 3-input AND.
 *
 *        X = ((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog wrapper for o221a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o221a_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o221a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O221A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o221ai: 2-input OR into first two inputs of 3-input NAND.
 *
 *         Y = !((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o221ai: 2-input OR into first two inputs of 3-input NAND.
 *
 *         Y = !((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o221ai (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire or1_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , B2, B1                 );
    or                                 or1         (or1_out          , A2, A1                 );
    nand                               nand0       (nand0_out_Y      , or1_out, or0_out, C1   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O221AI_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL



















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O221AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o221ai: 2-input OR into first two inputs of 3-input NAND.
 *
 *         Y = !((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog wrapper for o221ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o221ai_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o221ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O221AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o221ai: 2-input OR into first two inputs of 3-input NAND.
 *
 *         Y = !((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog wrapper for o221ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o221ai_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o221ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O221AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o221ai: 2-input OR into first two inputs of 3-input NAND.
 *
 *         Y = !((A1 | A2) & (B1 | B2) & C1)
 *
 * Verilog wrapper for o221ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o221ai_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o221ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O221AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311a: 3-input OR into 3-input AND.
 *
 *        X = ((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o311a: 3-input OR into 3-input AND.
 *
 *        X = ((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o311a (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1, A3            );
    and                                and0        (and0_out_X       , or0_out, B1, C1       );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O311A_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311a: 3-input OR into 3-input AND.
 *
 *        X = ((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog wrapper for o311a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o311a_1 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o311a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311a: 3-input OR into 3-input AND.
 *
 *        X = ((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog wrapper for o311a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o311a_2 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o311a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311a: 3-input OR into 3-input AND.
 *
 *        X = ((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog wrapper for o311a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o311a_4 (
    X   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o311a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311ai: 3-input OR into 3-input NAND.
 *
 *         Y = !((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o311ai: 3-input OR into 3-input NAND.
 *
 *         Y = !((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o311ai (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1, A3             );
    nand                               nand0       (nand0_out_Y      , C1, or0_out, B1        );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O311AI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311ai: 3-input OR into 3-input NAND.
 *
 *         Y = !((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog wrapper for o311ai with size of 0 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o311ai_0 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o311ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311AI_0_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311ai: 3-input OR into 3-input NAND.
 *
 *         Y = !((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog wrapper for o311ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o311ai_1 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o311ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311ai: 3-input OR into 3-input NAND.
 *
 *         Y = !((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog wrapper for o311ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o311ai_2 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o311ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o311ai: 3-input OR into 3-input NAND.
 *
 *         Y = !((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog wrapper for o311ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o311ai_4 (
    Y   ,
    A1  ,
    A2  ,
    A3  ,
    B1  ,
    C1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  B1  ;
    input  C1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o311ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .B1(B1),
        .C1(C1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O311AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2111a: 2-input OR into first input of 4-input AND.
 *
 *         X = ((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o2111a: 2-input OR into first input of 4-input AND.
 *
 *         X = ((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o2111a (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1                );
    and                                and0        (and0_out_X       , B1, C1, or0_out, D1   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O2111A_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2111A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2111a: 2-input OR into first input of 4-input AND.
 *
 *         X = ((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog wrapper for o2111a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2111a_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2111a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2111A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2111a: 2-input OR into first input of 4-input AND.
 *
 *         X = ((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog wrapper for o2111a with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2111a_2 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2111a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2111A_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2111a: 2-input OR into first input of 4-input AND.
 *
 *         X = ((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog wrapper for o2111a with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2111a_4 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2111a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2111A_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2111ai: 2-input OR into first input of 4-input NAND.
 *
 *          Y = !((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o2111ai: 2-input OR into first input of 4-input NAND.
 *
 *          Y = !((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__o2111ai (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out          , A2, A1                 );
    nand                               nand0       (nand0_out_Y      , C1, B1, D1, or0_out    );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__O2111AI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2111AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2111ai: 2-input OR into first input of 4-input NAND.
 *
 *          Y = !((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog wrapper for o2111ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2111ai_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2111ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2111AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2111ai: 2-input OR into first input of 4-input NAND.
 *
 *          Y = !((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog wrapper for o2111ai with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2111ai_2 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2111ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2111AI_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o2111ai: 2-input OR into first input of 4-input NAND.
 *
 *          Y = !((A1 | A2) & B1 & C1 & D1)
 *
 * Verilog wrapper for o2111ai with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__o2111ai_4 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    C1  ,
    D1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  C1  ;
    input  D1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__o2111ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .C1(C1),
        .D1(D1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__O2111AI_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2: 2-input OR.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or2: 2-input OR.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__or2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out_X        , B, A                 );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__OR2_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2: 2-input OR.
 *
 * Verilog wrapper for or2 with size of 0 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or2_0 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2_0_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2: 2-input OR.
 *
 * Verilog wrapper for or2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or2_1 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2: 2-input OR.
 *
 * Verilog wrapper for or2 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or2_2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2: 2-input OR.
 *
 * Verilog wrapper for or2 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or2_4 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2b: 2-input OR, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or2b: 2-input OR, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__or2b (
    X   ,
    A   ,
    B_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , B_N                  );
    or                                 or0         (or0_out_X        , not0_out, A          );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__OR2B_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2b: 2-input OR, first input inverted.
 *
 * Verilog wrapper for or2b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or2b_1 (
    X   ,
    A   ,
    B_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or2b base (
        .X(X),
        .A(A),
        .B_N(B_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2b: 2-input OR, first input inverted.
 *
 * Verilog wrapper for or2b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or2b_2 (
    X   ,
    A   ,
    B_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or2b base (
        .X(X),
        .A(A),
        .B_N(B_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2b: 2-input OR, first input inverted.
 *
 * Verilog wrapper for or2b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or2b_4 (
    X   ,
    A   ,
    B_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or2b base (
        .X(X),
        .A(A),
        .B_N(B_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR2B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3: 3-input OR.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or3: 3-input OR.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__or3 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out_X        , B, A, C              );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__OR3_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3: 3-input OR.
 *
 * Verilog wrapper for or3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or3_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3: 3-input OR.
 *
 * Verilog wrapper for or3 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or3_2 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR3_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3: 3-input OR.
 *
 * Verilog wrapper for or3 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or3_4 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR3_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3b: 3-input OR, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or3b: 3-input OR, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__or3b (
    X   ,
    A   ,
    B   ,
    C_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , C_N                  );
    or                                 or0         (or0_out_X        , B, A, not0_out       );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__OR3B_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR3B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3b: 3-input OR, first input inverted.
 *
 * Verilog wrapper for or3b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or3b_1 (
    X   ,
    A   ,
    B   ,
    C_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or3b base (
        .X(X),
        .A(A),
        .B(B),
        .C_N(C_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR3B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3b: 3-input OR, first input inverted.
 *
 * Verilog wrapper for or3b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or3b_2 (
    X   ,
    A   ,
    B   ,
    C_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or3b base (
        .X(X),
        .A(A),
        .B(B),
        .C_N(C_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR3B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3b: 3-input OR, first input inverted.
 *
 * Verilog wrapper for or3b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or3b_4 (
    X   ,
    A   ,
    B   ,
    C_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or3b base (
        .X(X),
        .A(A),
        .B(B),
        .C_N(C_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR3B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4: 4-input OR.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or4: 4-input OR.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__or4 (
    X   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    or                                 or0         (or0_out_X        , D, C, B, A           );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__OR4_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4: 4-input OR.
 *
 * Verilog wrapper for or4 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4: 4-input OR.
 *
 * Verilog wrapper for or4 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4_2 (
    X   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4: 4-input OR.
 *
 * Verilog wrapper for or4 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4_4 (
    X   ,
    A   ,
    B   ,
    C   ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4b: 4-input OR, first input inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or4b: 4-input OR, first input inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__or4b (
    X   ,
    A   ,
    B   ,
    C   ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    not                                not0        (not0_out         , D_N                  );
    or                                 or0         (or0_out_X        , not0_out, C, B, A    );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__OR4B_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4B_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4b: 4-input OR, first input inverted.
 *
 * Verilog wrapper for or4b with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4b_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4b base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4B_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4b: 4-input OR, first input inverted.
 *
 * Verilog wrapper for or4b with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4b_2 (
    X   ,
    A   ,
    B   ,
    C   ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4b base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4B_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4b: 4-input OR, first input inverted.
 *
 * Verilog wrapper for or4b with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4b_4 (
    X   ,
    A   ,
    B   ,
    C   ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4b base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4B_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4bb: 4-input OR, first two inputs inverted.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or4bb: 4-input OR, first two inputs inverted.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__or4bb (
    X   ,
    A   ,
    B   ,
    C_N ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    nand                               nand0       (nand0_out        , D_N, C_N             );
    or                                 or0         (or0_out_X        , B, A, nand0_out      );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__OR4BB_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4BB_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4bb: 4-input OR, first two inputs inverted.
 *
 * Verilog wrapper for or4bb with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4bb_1 (
    X   ,
    A   ,
    B   ,
    C_N ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4bb base (
        .X(X),
        .A(A),
        .B(B),
        .C_N(C_N),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4BB_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4bb: 4-input OR, first two inputs inverted.
 *
 * Verilog wrapper for or4bb with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4bb_2 (
    X   ,
    A   ,
    B   ,
    C_N ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4bb base (
        .X(X),
        .A(A),
        .B(B),
        .C_N(C_N),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4BB_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or4bb: 4-input OR, first two inputs inverted.
 *
 * Verilog wrapper for or4bb with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__or4bb_4 (
    X   ,
    A   ,
    B   ,
    C_N ,
    D_N ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C_N ;
    input  D_N ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__or4bb base (
        .X(X),
        .A(A),
        .B(B),
        .C_N(C_N),
        .D_N(D_N),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__OR4BB_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * probe_p: Virtual voltage probe point.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * probe_p: Virtual voltage probe point.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__probe_p (
    X   ,
    A   ,
    VGND,
    VNB ,
    VPB ,
    VPWR
);

    // Module ports
    output X   ;
    input  A   ;
    input  VGND;
    input  VNB ;
    input  VPB ;
    input  VPWR;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__PROBE_P_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__PROBE_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * probe_p: Virtual voltage probe point.
 *
 * Verilog wrapper for probe_p with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__probe_p_8 (
    X   ,
    A   ,
    VGND,
    VNB ,
    VPB ,
    VPWR
);

    output X   ;
    input  A   ;
    input  VGND;
    input  VNB ;
    input  VPB ;
    input  VPWR;
    sky130_fd_sc_hd__probe_p base (
        .X(X),
        .A(A),
        .VGND(VGND),
        .VNB(VNB),
        .VPB(VPB),
        .VPWR(VPWR)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__PROBE_P_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * probec_p: Virtual current probe point.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * probec_p: Virtual current probe point.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__probec_p (
    X   ,
    A   ,
    VGND,
    VNB ,
    VPB ,
    VPWR
);

    // Module ports
    output X   ;
    input  A   ;
    input  VGND;
    input  VNB ;
    input  VPB ;
    input  VPWR;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    buf                                buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__PROBEC_P_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__PROBEC_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * probec_p: Virtual current probe point.
 *
 * Verilog wrapper for probec_p with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__probec_p_8 (
    X   ,
    A   ,
    VGND,
    VNB ,
    VPB ,
    VPWR
);

    output X   ;
    input  A   ;
    input  VGND;
    input  VNB ;
    input  VPB ;
    input  VPWR;
    sky130_fd_sc_hd__probec_p base (
        .X(X),
        .A(A),
        .VGND(VGND),
        .VNB(VNB),
        .VPB(VPB),
        .VPWR(VPWR)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__PROBEC_P_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfbbn: Scan delay flop, inverted set, inverted reset, inverted
 *         clock, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfbbn: Scan delay flop, inverted set, inverted reset, inverted
 *         clock, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfbbn (
    Q      ,
    Q_N    ,
    D      ,
    SCD    ,
    SCE    ,
    CLK_N  ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  CLK_N  ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET  ;
    wire SET    ;
    wire CLK    ;
    wire buf_Q  ;
    wire mux_out;

    //                                   Delay       Name       Output   Other arguments
    not                                              not0      (RESET  , RESET_B                               );
    not                                              not1      (SET    , SET_B                                 );
    not                                              not2      (CLK    , CLK_N                                 );
    sky130_fd_sc_hd__udp_mux_2to1                    mux_2to10 (mux_out, D, SCD, SCE                           );
    sky130_fd_sc_hd__udp_dff$NSR_pp$PG$N #1 dff0      (buf_Q  , SET, RESET, CLK, mux_out, , VPWR, VGND);
    buf                                              buf0      (Q      , buf_Q                                 );
    not                                              not3      (Q_N    , buf_Q                                 );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFBBN_FUNCTIONAL_PP_V











































































































 // FUNCTIONAL




























































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFBBN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfbbn: Scan delay flop, inverted set, inverted reset, inverted
 *         clock, complementary outputs.
 *
 * Verilog wrapper for sdfbbn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfbbn_1 (
    Q      ,
    Q_N    ,
    D      ,
    SCD    ,
    SCE    ,
    CLK_N  ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  CLK_N  ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfbbn base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .CLK_N(CLK_N),
        .SET_B(SET_B),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/













































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFBBN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfbbn: Scan delay flop, inverted set, inverted reset, inverted
 *         clock, complementary outputs.
 *
 * Verilog wrapper for sdfbbn with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfbbn_2 (
    Q      ,
    Q_N    ,
    D      ,
    SCD    ,
    SCE    ,
    CLK_N  ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  CLK_N  ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfbbn base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .CLK_N(CLK_N),
        .SET_B(SET_B),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/













































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFBBN_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfbbp: Scan delay flop, inverted set, inverted reset, non-inverted
 *         clock, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfbbp: Scan delay flop, inverted set, inverted reset, non-inverted
 *         clock, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfbbp (
    Q      ,
    Q_N    ,
    D      ,
    SCD    ,
    SCE    ,
    CLK    ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  CLK    ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET  ;
    wire SET    ;
    wire buf_Q  ;
    wire mux_out;

    //                                   Delay       Name       Output   Other arguments
    not                                              not0      (RESET  , RESET_B                               );
    not                                              not1      (SET    , SET_B                                 );
    sky130_fd_sc_hd__udp_mux_2to1                    mux_2to10 (mux_out, D, SCD, SCE                           );
    sky130_fd_sc_hd__udp_dff$NSR_pp$PG$N #1 dff0      (buf_Q  , SET, RESET, CLK, mux_out, , VPWR, VGND);
    buf                                              buf0      (Q      , buf_Q                                 );
    not                                              not2      (Q_N    , buf_Q                                 );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFBBP_FUNCTIONAL_PP_V









































































































 // FUNCTIONAL
























































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFBBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfbbp: Scan delay flop, inverted set, inverted reset, non-inverted
 *         clock, complementary outputs.
 *
 * Verilog wrapper for sdfbbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfbbp_1 (
    Q      ,
    Q_N    ,
    D      ,
    SCD    ,
    SCE    ,
    CLK    ,
    SET_B  ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  CLK    ;
    input  SET_B  ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfbbp base (
        .Q(Q),
        .Q_N(Q_N),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .CLK(CLK),
        .SET_B(SET_B),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/













































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFBBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrbp: Scan delay flop, inverted reset, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfrbp: Scan delay flop, inverted reset, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfrbp (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q  ;
    wire RESET  ;
    wire mux_out;

    //                                  Delay       Name       Output   Other arguments
    not                                             not0      (RESET  , RESET_B                          );
    sky130_fd_sc_hd__udp_mux_2to1                   mux_2to10 (mux_out, D, SCD, SCE                      );
    sky130_fd_sc_hd__udp_dff$PR_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, RESET, , VPWR, VGND);
    buf                                             buf0      (Q      , buf_Q                            );
    not                                             not1      (Q_N    , buf_Q                            );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRBP_FUNCTIONAL_PP_V


































































































 // FUNCTIONAL













































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrbp: Scan delay flop, inverted reset, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog wrapper for sdfrbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfrbp_1 (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfrbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrbp: Scan delay flop, inverted reset, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog wrapper for sdfrbp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfrbp_2 (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfrbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRBP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrtn: Scan delay flop, inverted reset, inverted clock,
 *         single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfrtn: Scan delay flop, inverted reset, inverted clock,
 *         single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfrtn (
    Q      ,
    CLK_N  ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  CLK_N  ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q  ;
    wire RESET  ;
    wire intclk ;
    wire mux_out;

    //                                  Delay       Name       Output   Other arguments
    not                                             not0      (RESET  , RESET_B                             );
    not                                             not1      (intclk , CLK_N                               );
    sky130_fd_sc_hd__udp_mux_2to1                   mux_2to10 (mux_out, D, SCD, SCE                         );
    sky130_fd_sc_hd__udp_dff$PR_pp$PG$N #1 dff0      (buf_Q  , mux_out, intclk, RESET, , VPWR, VGND);
    buf                                             buf0      (Q      , buf_Q                               );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRTN_FUNCTIONAL_PP_V

































































































 // FUNCTIONAL











































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRTN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrtn: Scan delay flop, inverted reset, inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfrtn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfrtn_1 (
    Q      ,
    CLK_N  ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK_N  ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfrtn base (
        .Q(Q),
        .CLK_N(CLK_N),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRTN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrtp: Scan delay flop, inverted reset, non-inverted clock,
 *         single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfrtp: Scan delay flop, inverted reset, non-inverted clock,
 *         single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfrtp (
    Q      ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q  ;
    wire RESET  ;
    wire mux_out;

    //                                  Delay       Name       Output   Other arguments
    not                                             not0      (RESET  , RESET_B                          );
    sky130_fd_sc_hd__udp_mux_2to1                   mux_2to10 (mux_out, D, SCD, SCE                      );
    sky130_fd_sc_hd__udp_dff$PR_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, RESET, , VPWR, VGND);
    buf                                             buf0      (Q      , buf_Q                            );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRTP_FUNCTIONAL_PP_V































































































 // FUNCTIONAL







































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrtp: Scan delay flop, inverted reset, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfrtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfrtp_1 (
    Q      ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfrtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrtp: Scan delay flop, inverted reset, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfrtp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfrtp_2 (
    Q      ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfrtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRTP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrtp: Scan delay flop, inverted reset, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfrtp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfrtp_4 (
    Q      ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hd__sdfrtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFRTP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfsbp: Scan delay flop, inverted set, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfsbp: Scan delay flop, inverted set, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfsbp (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf_Q  ;
    wire SET    ;
    wire mux_out;

    //                                  Delay       Name       Output   Other arguments
    not                                             not0      (SET    , SET_B                          );
    sky130_fd_sc_hd__udp_mux_2to1                   mux_2to10 (mux_out, D, SCD, SCE                    );
    sky130_fd_sc_hd__udp_dff$PS_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, SET, , VPWR, VGND);
    buf                                             buf0      (Q      , buf_Q                          );
    not                                             not1      (Q_N    , buf_Q                          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSBP_FUNCTIONAL_PP_V


































































































 // FUNCTIONAL













































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfsbp: Scan delay flop, inverted set, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog wrapper for sdfsbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfsbp_1 (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__sdfsbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfsbp: Scan delay flop, inverted set, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog wrapper for sdfsbp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfsbp_2 (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__sdfsbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSBP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfstp: Scan delay flop, inverted set, non-inverted clock,
 *         single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfstp: Scan delay flop, inverted set, non-inverted clock,
 *         single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfstp (
    Q    ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf_Q  ;
    wire SET    ;
    wire mux_out;

    //                                  Delay       Name       Output   Other arguments
    not                                             not0      (SET    , SET_B                          );
    sky130_fd_sc_hd__udp_mux_2to1                   mux_2to10 (mux_out, D, SCD, SCE                    );
    sky130_fd_sc_hd__udp_dff$PS_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, SET, , VPWR, VGND);
    buf                                             buf0      (Q      , buf_Q                          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSTP_FUNCTIONAL_PP_V































































































 // FUNCTIONAL







































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfstp: Scan delay flop, inverted set, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfstp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfstp_1 (
    Q    ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__sdfstp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfstp: Scan delay flop, inverted set, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfstp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfstp_2 (
    Q    ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__sdfstp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSTP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfstp: Scan delay flop, inverted set, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfstp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfstp_4 (
    Q    ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hd__sdfstp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFSTP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxbp: Scan delay flop, non-inverted clock, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfxbp: Scan delay flop, non-inverted clock, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfxbp (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q  ;
    wire mux_out;

    //                                 Delay       Name       Output   Other arguments
    sky130_fd_sc_hd__udp_mux_2to1                  mux_2to10 (mux_out, D, SCD, SCE               );
    sky130_fd_sc_hd__udp_dff$P_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, , VPWR, VGND);
    buf                                            buf0      (Q      , buf_Q                     );
    not                                            not0      (Q_N    , buf_Q                     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXBP_FUNCTIONAL_PP_V
























































































 // FUNCTIONAL






























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxbp: Scan delay flop, non-inverted clock, complementary outputs.
 *
 * Verilog wrapper for sdfxbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfxbp_1 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sdfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxbp: Scan delay flop, non-inverted clock, complementary outputs.
 *
 * Verilog wrapper for sdfxbp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfxbp_2 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sdfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXBP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxtp: Scan delay flop, non-inverted clock, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfxtp: Scan delay flop, non-inverted clock, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdfxtp (
    Q   ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q  ;
    wire mux_out;

    //                                 Delay       Name       Output   Other arguments
    sky130_fd_sc_hd__udp_mux_2to1                  mux_2to10 (mux_out, D, SCD, SCE               );
    sky130_fd_sc_hd__udp_dff$P_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, , VPWR, VGND);
    buf                                            buf0      (Q      , buf_Q                     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXTP_FUNCTIONAL_PP_V





















































































 // FUNCTIONAL
























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxtp: Scan delay flop, non-inverted clock, single output.
 *
 * Verilog wrapper for sdfxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfxtp_1 (
    Q   ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sdfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxtp: Scan delay flop, non-inverted clock, single output.
 *
 * Verilog wrapper for sdfxtp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfxtp_2 (
    Q   ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sdfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXTP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxtp: Scan delay flop, non-inverted clock, single output.
 *
 * Verilog wrapper for sdfxtp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdfxtp_4 (
    Q   ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sdfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDFXTP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdlclkp: Scan gated clock.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdlclkp: Scan gated clock.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sdlclkp (
    GCLK,
    SCE ,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output GCLK;
    input  SCE ;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire m0      ;
    wire m0n     ;
    wire clkn    ;
    wire SCE_GATE;

    //                                    Name     Output    Other arguments
    not                                   not0    (m0n     , m0                          );
    not                                   not1    (clkn    , CLK                         );
    nor                                   nor0    (SCE_GATE, GATE, SCE                   );
    sky130_fd_sc_hd__udp_dlatch$P_pp$PG$N dlatch0 (m0      , SCE_GATE, clkn, , VPWR, VGND);
    and                                   and0    (GCLK    , m0n, CLK                    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SDLCLKP_FUNCTIONAL_PP_V




















































































 // FUNCTIONAL

























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDLCLKP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdlclkp: Scan gated clock.
 *
 * Verilog wrapper for sdlclkp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdlclkp_1 (
    GCLK,
    SCE ,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output GCLK;
    input  SCE ;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sdlclkp base (
        .GCLK(GCLK),
        .SCE(SCE),
        .GATE(GATE),
        .CLK(CLK),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDLCLKP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdlclkp: Scan gated clock.
 *
 * Verilog wrapper for sdlclkp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdlclkp_2 (
    GCLK,
    SCE ,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output GCLK;
    input  SCE ;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sdlclkp base (
        .GCLK(GCLK),
        .SCE(SCE),
        .GATE(GATE),
        .CLK(CLK),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDLCLKP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdlclkp: Scan gated clock.
 *
 * Verilog wrapper for sdlclkp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sdlclkp_4 (
    GCLK,
    SCE ,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output GCLK;
    input  SCE ;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sdlclkp base (
        .GCLK(GCLK),
        .SCE(SCE),
        .GATE(GATE),
        .CLK(CLK),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SDLCLKP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sedfxbp: Scan delay flop, data enable, non-inverted clock,
 *          complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sedfxbp: Scan delay flop, data enable, non-inverted clock,
 *          complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sedfxbp (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    DE  ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q  ;
    wire mux_out;
    wire de_d   ;

    //                                 Delay       Name       Output   Other arguments
    sky130_fd_sc_hd__udp_mux_2to1                  mux_2to10 (mux_out, de_d, SCD, SCE            );
    sky130_fd_sc_hd__udp_mux_2to1                  mux_2to11 (de_d   , buf_Q, D, DE              );
    sky130_fd_sc_hd__udp_dff$P_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, , VPWR, VGND);
    buf                                            buf0      (Q      , buf_Q                     );
    not                                            not0      (Q_N    , buf_Q                     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXBP_FUNCTIONAL_PP_V






























































































 // FUNCTIONAL









































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sedfxbp: Scan delay flop, data enable, non-inverted clock,
 *          complementary outputs.
 *
 * Verilog wrapper for sedfxbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sedfxbp_1 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    DE  ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sedfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .DE(DE),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sedfxbp: Scan delay flop, data enable, non-inverted clock,
 *          complementary outputs.
 *
 * Verilog wrapper for sedfxbp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sedfxbp_2 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    DE  ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sedfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .DE(DE),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXBP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sedfxtp: Scan delay flop, data enable, non-inverted clock,
 *          single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sedfxtp: Scan delay flop, data enable, non-inverted clock,
 *          single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__sedfxtp (
    Q   ,
    CLK ,
    D   ,
    DE  ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q  ;
    wire mux_out;
    wire de_d   ;

    //                                 Delay       Name       Output   Other arguments
    sky130_fd_sc_hd__udp_mux_2to1                  mux_2to10 (mux_out, de_d, SCD, SCE            );
    sky130_fd_sc_hd__udp_mux_2to1                  mux_2to11 (de_d   , buf_Q, D, DE              );
    sky130_fd_sc_hd__udp_dff$P_pp$PG$N #1 dff0      (buf_Q  , mux_out, CLK, , VPWR, VGND);
    buf                                            buf0      (Q      , buf_Q                     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXTP_FUNCTIONAL_PP_V



























































































 // FUNCTIONAL



































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sedfxtp: Scan delay flop, data enable, non-inverted clock,
 *          single output.
 *
 * Verilog wrapper for sedfxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sedfxtp_1 (
    Q   ,
    CLK ,
    D   ,
    DE  ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sedfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .DE(DE),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sedfxtp: Scan delay flop, data enable, non-inverted clock,
 *          single output.
 *
 * Verilog wrapper for sedfxtp with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sedfxtp_2 (
    Q   ,
    CLK ,
    D   ,
    DE  ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sedfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .DE(DE),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXTP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sedfxtp: Scan delay flop, data enable, non-inverted clock,
 *          single output.
 *
 * Verilog wrapper for sedfxtp with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__sedfxtp_4 (
    Q   ,
    CLK ,
    D   ,
    DE  ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  DE  ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__sedfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .DE(DE),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__SEDFXTP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tap: Tap cell with no tap connections (no contacts on metal1).
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * tap: Tap cell with no tap connections (no contacts on metal1).
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__tap (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__TAP_FUNCTIONAL_PP_V



















































 // FUNCTIONAL



























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tap: Tap cell with no tap connections (no contacts on metal1).
 *
 * Verilog wrapper for tap with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__tap_1 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__tap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tap: Tap cell with no tap connections (no contacts on metal1).
 *
 * Verilog wrapper for tap with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__tap_2 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__tap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAP_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tapvgnd2: Tap cell with tap to ground, isolated power connection
 *           2 rows down.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * tapvgnd2: Tap cell with tap to ground, isolated power connection 2
 *           rows down.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__tapvgnd2 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVGND2_FUNCTIONAL_PP_V




















































 // FUNCTIONAL





























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVGND2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tapvgnd2: Tap cell with tap to ground, isolated power connection
 *           2 rows down.
 *
 * Verilog wrapper for tapvgnd2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__tapvgnd2_1 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__tapvgnd2 base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVGND2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tapvgnd: Tap cell with tap to ground, isolated power connection
 *          1 row down.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * tapvgnd: Tap cell with tap to ground, isolated power connection 1
 *          row down.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__tapvgnd (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVGND_FUNCTIONAL_PP_V




















































 // FUNCTIONAL





























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVGND_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tapvgnd: Tap cell with tap to ground, isolated power connection
 *          1 row down.
 *
 * Verilog wrapper for tapvgnd with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__tapvgnd_1 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__tapvgnd base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVGND_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tapvpwrvgnd: Substrate and well tap cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * tapvpwrvgnd: Substrate and well tap cell.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hd__tapvpwrvgnd (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVPWRVGND_FUNCTIONAL_PP_V



















































 // FUNCTIONAL



























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVPWRVGND_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * tapvpwrvgnd: Substrate and well tap cell.
 *
 * Verilog wrapper for tapvpwrvgnd with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__tapvpwrvgnd_1 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hd__tapvpwrvgnd base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__TAPVPWRVGND_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor2: 2-input exclusive NOR.
 *
 *        Y = !(A ^ B)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * xnor2: 2-input exclusive NOR.
 *
 *        Y = !(A ^ B)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__xnor2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire xnor0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                 Name         Output             Other arguments
    xnor                               xnor0       (xnor0_out_Y      , A, B                   );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, xnor0_out_Y, VPWR, VGND);
    buf                                buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR2_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor2: 2-input exclusive NOR.
 *
 *        Y = !(A ^ B)
 *
 * Verilog wrapper for xnor2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xnor2_1 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xnor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor2: 2-input exclusive NOR.
 *
 *        Y = !(A ^ B)
 *
 * Verilog wrapper for xnor2 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xnor2_2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xnor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR2_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor2: 2-input exclusive NOR.
 *
 *        Y = !(A ^ B)
 *
 * Verilog wrapper for xnor2 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xnor2_4 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xnor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR2_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor3: 3-input exclusive NOR.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * xnor3: 3-input exclusive NOR.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__xnor3 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire xnor0_out_X      ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    xnor                               xnor0       (xnor0_out_X      , A, B, C                );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, xnor0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR3_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor3: 3-input exclusive NOR.
 *
 * Verilog wrapper for xnor3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xnor3_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xnor3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor3: 3-input exclusive NOR.
 *
 * Verilog wrapper for xnor3 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xnor3_2 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xnor3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR3_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor3: 3-input exclusive NOR.
 *
 * Verilog wrapper for xnor3 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xnor3_4 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xnor3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XNOR3_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor2: 2-input exclusive OR.
 *
 *       X = A ^ B
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * xor2: 2-input exclusive OR.
 *
 *       X = A ^ B
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__xor2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire xor0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    xor                                xor0        (xor0_out_X       , B, A                  );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, xor0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__XOR2_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XOR2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor2: 2-input exclusive OR.
 *
 *       X = A ^ B
 *
 * Verilog wrapper for xor2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xor2_1 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xor2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XOR2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor2: 2-input exclusive OR.
 *
 *       X = A ^ B
 *
 * Verilog wrapper for xor2 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xor2_2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xor2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XOR2_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor2: 2-input exclusive OR.
 *
 *       X = A ^ B
 *
 * Verilog wrapper for xor2 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xor2_4 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xor2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XOR2_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor3: 3-input exclusive OR.
 *
 *       X = A ^ B ^ C
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * xor3: 3-input exclusive OR.
 *
 *       X = A ^ B ^ C
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hd__xor3 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire xor0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                 Name         Output             Other arguments
    xor                                xor0        (xor0_out_X       , A, B, C               );
    sky130_fd_sc_hd__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, xor0_out_X, VPWR, VGND);
    buf                                buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HD__XOR3_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XOR3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor3: 3-input exclusive OR.
 *
 *       X = A ^ B ^ C
 *
 * Verilog wrapper for xor3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xor3_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xor3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XOR3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor3: 3-input exclusive OR.
 *
 *       X = A ^ B ^ C
 *
 * Verilog wrapper for xor3 with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xor3_2 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xor3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XOR3_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor3: 3-input exclusive OR.
 *
 *       X = A ^ B ^ C
 *
 * Verilog wrapper for xor3 with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hd__xor3_4 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hd__xor3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HD__XOR3_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$P: Positive edge triggered D flip-flop (Q output UDP).
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dff$P (
    Q  ,
    D  ,
    CLK
);

    output Q  ;
    input  D  ;
    input  CLK;

    reg Q;

    table
     //  D  CLK  :  Qt : Qt+1
         1  (01) :  ?  :  1    ; // clocked data
         0  (01) :  ?  :  0    ;
         1  (x1) :  1  :  1    ; // reducing pessimism
         0  (x1) :  0  :  0    ;
         0   x   :  0  :  0    ; // unkown CP, hold when D==Q==0
         1   x   :  1  :  1    ; // unkown CP, hold when D==Q==1
         ?  (?0) :  ?  :  -    ;
         *   b   :  ?  :  -    ; // ignore edges on data, unless CP=X
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DFF_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$P_pp$PG$N: Positive edge triggered D flip-flop
 *                    (Q output UDP).
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dff$P_pp$PG$N (
    Q       ,
    D       ,
    CLK     ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  CLK     ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           CLK  NOTIFIER VPWR VGND :  Qt : Qt+1
                 1           (01)    ?      1    0   :  ?  :  1    ; // clocked data
                 0           (01)    ?      1    0   :  ?  :  0    ;
                 1           (x1)    ?      1    0   :  1  :  1    ; // reducing pessimism
                 0           (x1)    ?      1    0   :  0  :  0    ;
                 1           (0x)    ?      1    0   :  1  :  1    ;
                 0           (0x)    ?      1    0   :  0  :  0    ;
                 0            x      ?      1    0   :  0  :  0    ; // Hold when CLK=X and D=Q
                 1            x      ?      1    0   :  1  :  1    ; // Hold when CLK=X and D=Q
                 ?           (?0)    ?      1    0   :  ?  :  -    ;
                 *            b      ?      1    0   :  ?  :  -    ; // ignore edges on data
        // ['IfDef(functional)', '']                 ?            ?      *      1    0   :  ?  :  -    ;
        // ['Else', '']                 ?            ?      *      1    0   :  ?  :  x    ;
        // ['EndIfDef(functional)', '']                 ?            ?      ?      *    ?   :  ?  :  x    ; // any change on vpwr
                 ?            ?      ?      ?    *   :  ?  :  x    ; // any change on vgnd
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DFF_P_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$PR: Positive edge triggered D flip-flop with active high
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dff$PR (
    Q    ,
    D    ,
    CLK  ,
    RESET
);

    output Q    ;
    input  D    ;
    input  CLK  ;
    input  RESET;

    reg Q;

    table
     //  D  CLK  RESET :  Qt : Qt+1
         *   b     0   :  ?  :  -    ; // data event, hold unless CP==x
         ?  (?0)   0   :  ?  :  -    ; // CP => 0, hold
         ?   b    (?0) :  ?  :  -    ; // R => 0, hold unless CP==x
         ?   ?     1   :  ?  :  0    ; // async reset
         0   r     ?   :  ?  :  0    ; // clock data on CP
         1   r     0   :  ?  :  1    ; // clock data on CP
         0  (x1)   ?   :  0  :  0    ; // possible CP, hold when D==Q==0
         1  (x1)   0   :  1  :  1    ; // possible CP, hold when D==Q==1
         0   x     ?   :  0  :  0    ; // unkown CP, hold when D==Q==0
         1   x     0   :  1  :  1    ; // unkown CP, hold when D==Q==1
         ?   b    (?x) :  0  :  0    ; // R=>x, hold when Q==0 unless CP==x
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DFF_PR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$PR_pp$PG$N: Positive edge triggered D flip-flop with active
 *                     high
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dff$PR_pp$PG$N (
    Q       ,
    D       ,
    CLK     ,
    RESET   ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  CLK     ;
    input  RESET   ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           CLK  RESET NOTIFIER VPWR VGND :  Qt : Qt+1
                 *            b     0      ?      1    0   :  ?  :  -    ; // data event, hold unless CP==x
                 ?           (?0)   0      ?      1    0   :  ?  :  -    ; // CP => 0, hold
                 ?            b    (?0)    ?      1    0   :  ?  :  -    ; // R => 0, hold unless CP==x
                 ?            ?     1      ?      1    0   :  ?  :  0    ; // async reset
                 0            r     ?      ?      1    0   :  ?  :  0    ; // clock data on CP
                 1            r     0      ?      1    0   :  ?  :  1    ; // clock data on CP
                 0           (x1)   ?      ?      1    0   :  0  :  0    ; // possible CP, hold when D==Q==0
                 1           (x1)   0      ?      1    0   :  1  :  1    ; // possible CP, hold when D==Q==1
                 0            x     ?      ?      1    0   :  0  :  0    ; // unkown CP, hold when D==Q==0
                 1            x     0      ?      1    0   :  1  :  1    ; // unkown CP, hold when D==Q==1
                 ?            b    (?x)    ?      1    0   :  0  :  0    ; // R=>x, hold when Q==0 unless CP==x
                 ?            f     x      ?      1    0   :  0  :  0    ; // JCWR reducing pessimism
        // ['IfDef(functional)', '']                 ?            ?     ?      *      1    0   :  ?  :  -    ; // ignore notifier
        // ['Else', '']                 ?            ?     ?      *      1    0   :  ?  :  x    ; // Q => X on any change on notifier
        // ['EndIfDef(functional)', '']                 ?            ?     ?      ?      *    ?   :  ?  :  x    ; // Q => X on any change on vpwr
                 ?            ?     ?      ?      ?    *   :  ?  :  x    ; // Q => X on any change on vgnd
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DFF_PR_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$PS: Positive edge triggered D flip-flop with active high
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dff$PS (
    Q  ,
    D  ,
    CLK,
    SET
);

    output Q  ;
    input  D  ;
    input  CLK;
    input  SET;

    reg Q;

    table
     //  D  CLK  SET  :  Qt : Qt+1
         *   b    0   :  ?  :  -    ; // data event, hold unless CP==x
         ?  (?0)  0   :  ?  :  -    ; // CP => 0, hold
         ?   b   (?0) :  ?  :  -    ; // S => 0, hold unless CP==x
         ?   ?    1   :  ?  :  1    ; // async set
         0   r    0   :  ?  :  0    ; // clock data on CP
         1   r    ?   :  ?  :  1    ; // clock data on CP
         0  (x1)  0   :  0  :  0    ; // possible CP, hold when D==Q==0
         1  (x1)  ?   :  1  :  1    ; // possible CP, hold when D==Q==1
         0   x    0   :  0  :  0    ; // unkown CP, hold when D==Q==0
         1   x    ?   :  1  :  1    ; // unkown CP, hold when D==Q==1
         ?   b   (?x) :  1  :  1    ; // S=>x, hold when Q==1 unless CP==x
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DFF_PS_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dff$PS_pp$PG$N: Positive edge triggered D flip-flop with active
 *                     high
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dff$PS_pp$PG$N (
    Q       ,
    D       ,
    CLK     ,
    SET     ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  CLK     ;
    input  SET     ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           CLK  SET  NOTIFIER VPWR VGND :  Qt : Qt+1
                 *            b    0      ?      1    0   :  ?  :  -    ; // data event, hold unless CP==x
                 ?           (?0)  0      ?      1    0   :  ?  :  -    ; // CP => 0, hold
                 ?            b   (?0)    ?      1    0   :  ?  :  -    ; // S => 0, hold unless CP==x
                 ?            ?    1      ?      1    0   :  ?  :  1    ; // async set
                 0            r    0      ?      1    0   :  ?  :  0    ; // clock data on CP
                 1            r    ?      ?      1    0   :  ?  :  1    ; // clock data on CP
                 0           (x1)  0      ?      1    0   :  0  :  0    ; // possible CP, hold when D==Q==0
                 1           (x1)  ?      ?      1    0   :  1  :  1    ; // possible CP, hold when D==Q==1
                 0            x    0      ?      1    0   :  0  :  0    ; // unkown CP, hold when D==Q==0
                 1            x    ?      ?      1    0   :  1  :  1    ; // unkown CP, hold when D==Q==1
                 ?            b   (?x)    ?      1    0   :  1  :  1    ; // S=>x, hold when Q==1 unless CP==x
                 ?            f    x      ?      1    0   :  1  :  1    ; // JCWR reducing pessimism
        // ['IfDef(functional)', '']                 ?            ?    ?      *      1    0   :  ?  :  -    ; // ignore notifier
        // ['Else', '']                 ?            ?    ?      *      1    0   :  ?  :  x    ; // Q => X on any change on notifier
        // ['EndIfDef(functional)', '']                 ?            ?    ?      ?      *    ?   :  ?  :  x    ; // Q => X on any change on vpwr
                 ?            ?    ?      ?      ?    *   :  ?  :  x    ; // Q => X on any change on vgnd
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DFF_PS_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$P: D-latch, gated standard drive / active high
 *               (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dlatch$P (
    Q   ,
    D   ,
    GATE
);

    output Q   ;
    input  D   ;
    input  GATE;

    reg Q;

    table
     //  D  GATE :  Qt : Qt+1
         ?   0   :  ?  :  -    ; // hold
         0   1   :  ?  :  0    ; // pass 0
         1   1   :  ?  :  1    ; // pass 1
         0   x   :  0  :  0    ; // reduce pessimism
         1   x   :  1  :  1    ; // reduce pessimism
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DLATCH_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$P_pp$PG$N: D-latch, gated standard drive / active high
 *                       (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dlatch$P_pp$PG$N (
    Q       ,
    D       ,
    GATE    ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  GATE    ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           GATE NOTIFIER VPWR VGND : Qtn : Qtn+1
                 *            0      ?      1    0   :  ?  :   -    ;
                 ?           (?0)    ?      1    0   :  ?  :   -    ;
                 ?           (1x)    ?      1    0   :  ?  :   -    ;
                 0           (0x)    ?      1    0   :  0  :   0    ;
                 1           (0x)    ?      1    0   :  1  :   1    ;
                 0           (x1)    ?      1    0   :  ?  :   0    ;
                 1           (x1)    ?      1    0   :  ?  :   1    ;
                 0            1      ?      1    0   :  ?  :   0    ;
                 1            1      ?      1    0   :  ?  :   1    ;
                 0           (01)    ?      1    0   :  ?  :   0    ;
                 1           (01)    ?      1    0   :  ?  :   1    ;
                 1            x      ?      1    0   :  1  :   1    ; // Reducing pessimism.
                 0            x      ?      1    0   :  0  :   0    ;
        // ['IfDef(functional)', '']                 ?            ?      *      1    0   :  ?  :   -    ; // ignore notifier
        // ['Else', '']                 ?            ?      *      1    0   :  ?  :   x    ; // notifier
        // ['EndIfDef(functional)', '']                 ?            ?      ?      0    ?   :  ?  :   x    ; // vpwr != 1
                 ?            ?      ?      x    ?   :  ?  :   x    ; // vpwr != 1
                 ?            ?      ?      ?    1   :  ?  :   x    ; // vgnd != 0
                 ?            ?      ?      ?    x   :  ?  :   x    ; // vgnd != 0
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DLATCH_P_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$PR: D-latch, gated clear direct / gate active high
 *                (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dlatch$PR (
    Q    ,
    D    ,
    GATE ,
    RESET
);

    output Q    ;
    input  D    ;
    input  GATE ;
    input  RESET;

    reg Q;

    table
     //  D  GATE RESET :  Qt : Qt+1
         ?   0     0   :  ?  :  -    ; // hold
         0   1     0   :  ?  :  0    ; // pass 0
         1   1     0   :  ?  :  1    ; // pass 1
         ?   ?     1   :  ?  :  0    ; // async reset
         0   1     ?   :  ?  :  0    ; // reduce pessimism
         0   x     0   :  0  :  0    ; // reduce pessimism
         1   x     0   :  1  :  1    ; // reduce pessimism
         ?   0     x   :  0  :  0    ; // reduce pessimism
         0   x     x   :  0  :  0    ; // reduce pessimism
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DLATCH_PR_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_dlatch$PR_pp$PG$N: D-latch, gated clear direct / gate active
 *                        high (Q output UDP)
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_dlatch$PR_pp$PG$N (
    Q       ,
    D       ,
    GATE    ,
    RESET   ,
    NOTIFIER,
    VPWR    ,
    VGND
);

    output Q       ;
    input  D       ;
    input  GATE    ;
    input  RESET   ;
    input  NOTIFIER;
    input  VPWR    ;
    input  VGND    ;

    reg Q;

    table
     //          D           GATE RESET NOTIFIER VPWR VGND :  Qt : Qt+1
                 *            0     0      ?      1    0   :  ?  :  -    ;
                 ?            ?     1      ?      1    0   :  ?  :  0    ; // asynchro clear
                 ?           (?0)   0      ?      1    0   :  ?  :  -    ; // Changed R=? to R=0 ; jek 08/14/06/
                 ?           (1x)   0      ?      1    0   :  ?  :  -    ; // Changed R=? to R=0 ; jek 08/14/06
                 0           (0x)   0      ?      1    0   :  0  :  0    ;
                 1           (0x)   0      ?      1    0   :  1  :  1    ;
                 0           (x1)   0      ?      1    0   :  ?  :  0    ;
                 1           (x1)   0      ?      1    0   :  ?  :  1    ;
                 0            1     0      ?      1    0   :  ?  :  0    ;
                 1            1     0      ?      1    0   :  ?  :  1    ;
                 0           (01)   0      ?      1    0   :  ?  :  0    ;
                 1           (01)   0      ?      1    0   :  ?  :  1    ;
                 ?            0    (?x)    ?      1    0   :  0  :  0    ; // Reducing pessimism.//AB
                 *            0     x      ?      1    0   :  0  :  0    ; // Reducing pessimism//AB
                 0           (?1)   x      ?      1    0   :  ?  :  0    ; // Reducing pessimism.
                (?0)          1     x      ?      1    0   :  ?  :  0    ; // Reducing pessimism.
                 0            1    (?x)    ?      1    0   :  ?  :  0    ; // Reducing pessimism.//AB
                 ?            0    (?0)    ?      1    0   :  ?  :  -    ; // ignore edge on clear
                 0            1    (?0)    ?      1    0   :  ?  :  0    ; // pessimism .
                 1            1    (?0)    ?      1    0   :  ?  :  1    ;
                 1            x     0      ?      1    0   :  1  :  1    ; // Reducing pessimism.
                 0            x     0      ?      1    0   :  0  :  0    ; // Reducing pessimism.
        // ['IfDef(functional)', '']                 ?            ?     ?      *      1    0   :  ?  :  -    ; // ignore notifier
        // ['Else', '']                 ?            ?     ?      *      1    0   :  ?  :  x    ; // notifier
        // ['EndIfDef(functional)', '']                 ?            ?     ?      ?      0    ?   :  ?  :  x    ; // vpwr != 1
                 ?            ?     ?      ?      x    ?   :  ?  :  x    ; // vpwr != 1
                 ?            ?     ?      ?      ?    1   :  ?  :  x    ; // vgnd != 0
                 ?            ?     ?      ?      ?    x   :  ?  :  x    ; // vgnd != 0
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_DLATCH_PR_PP_PG_N_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_isolatchhv_pp$PLG$S: Power isolating latch (for HV). Includes
 *                          VPWR, LVPWR, and VGND power pins with
 *                          active high sleep pin (SLEEP).
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_isolatchhv_pp$PLG$S (
    UDP_OUT,
    UDP_IN ,
    VPWR   ,
    LVPWR  ,
    VGND   ,
    SLEEP
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VPWR   ;
    input  LVPWR  ;
    input  VGND   ;
    input  SLEEP  ;

    table
     // UDP_IN VPWR LVPWR VGND SLEEP : out
          0     1     1    0     b   :  0   ;
          1     1     1    0     0   :  1   ;
          b     1     ?    0     1   :  0   ;
          ?     1     0    0     1   :  0   ;
          x     1     1    0     1   :  x   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_ISOLATCHHV_PP_PLG_S_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_mux_2to1: Two to one multiplexer
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_mux_2to1 (
    X ,
    A0,
    A1,
    S
);

    output X ;
    input  A0;
    input  A1;
    input  S ;

    table
     //  A0  A1  S  :  X
         0   0   ?  :  0   ;
         1   1   ?  :  1   ;
         0   ?   0  :  0   ;
         1   ?   0  :  1   ;
         ?   0   1  :  0   ;
         ?   1   1  :  1   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_MUX_2TO1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * udp_mux_4to2: Four to one multiplexer with 2 select controls
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_mux_4to2 (
    X ,
    A0,
    A1,
    A2,
    A3,
    S0,
    S1
);

    output X ;
    input  A0;
    input  A1;
    input  A2;
    input  A3;
    input  S0;
    input  S1;

    table
     //  A0  A1  A2  A3  S0  S1 :  X
         0   ?   ?   ?   0   0  :  0   ;
         1   ?   ?   ?   0   0  :  1   ;
         ?   0   ?   ?   1   0  :  0   ;
         ?   1   ?   ?   1   0  :  1   ;
         ?   ?   0   ?   0   1  :  0   ;
         ?   ?   1   ?   0   1  :  1   ;
         ?   ?   ?   0   1   1  :  0   ;
         ?   ?   ?   1   1   1  :  1   ;
         0   0   0   0   ?   ?  :  0   ;
         1   1   1   1   ?   ?  :  1   ;
         0   0   ?   ?   ?   0  :  0   ;
         1   1   ?   ?   ?   0  :  1   ;
         ?   ?   0   0   ?   1  :  0   ;
         ?   ?   1   1   ?   1  :  1   ;
         0   ?   0   ?   0   ?  :  0   ;
         1   ?   1   ?   0   ?  :  1   ;
         ?   0   ?   0   1   ?  :  0   ;
         ?   1   ?   1   1   ?  :  1   ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_MUX_4TO2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VPWR!=1
 *   UDP_OUT :=UDP_IN when VPWR==1
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_pwrgood_pp$G (
    UDP_OUT,
    UDP_IN ,
    VGND
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VGND   ;

    table
     // UDP_IN VPWR : UDP_OUT
          0     0   :    0     ;
          1     0   :    1     ;
          ?     1   :    x     ;
          ?     x   :    x     ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_PWRGOOD_PP_G_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VPWR!=1
 *   UDP_OUT :=UDP_IN when VPWR==1
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_pwrgood_pp$P (
    UDP_OUT,
    UDP_IN ,
    VPWR
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VPWR   ;

    table
     // UDP_IN VPWR : UDP_OUT
          0     1   :    0     ;
          1     1   :    1     ;
          ?     0   :    x     ;
          ?     x   :    x     ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_PWRGOOD_PP_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**

 *   UDP_OUT :=x when VPWR!=1 or VGND!=0
 *   UDP_OUT :=UDP_IN when VPWR==1 and VGND==0
 *
 * Verilog primitive definition.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



primitive sky130_fd_sc_hvl__udp_pwrgood_pp$PG (
    UDP_OUT,
    UDP_IN ,
    VPWR   ,
    VGND
);

    output UDP_OUT;
    input  UDP_IN ;
    input  VPWR   ;
    input  VGND   ;

    table
     // UDP_IN VPWR VGND : UDP_OUT
          0     1    0   :    0     ;
          1     1    0   :    1     ;
          1     0    0   :    x     ;
          1     1    1   :    x     ;
          1     x    0   :    x     ;
          1     1    x   :    x     ;
    endtable
endprimitive
 // NO_PRIMITIVES

`default_nettype wire
  // SKY130_FD_SC_HVL__UDP_PWRGOOD_PP_PG_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21o: 2-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2) | B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a21o: 2-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2) | B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__a21o (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    and                                 and0        (and0_out         , A1, A2               );
    or                                  or0         (or0_out_X        , and0_out, B1         );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__A21O_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__A21O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21o: 2-input AND into first input of 2-input OR.
 *
 *       X = ((A1 & A2) | B1)
 *
 * Verilog wrapper for a21o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__a21o_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__a21o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__A21O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21oi: 2-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2) | B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a21oi: 2-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2) | B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__a21oi (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    and                                 and0        (and0_out         , A1, A2                );
    nor                                 nor0        (nor0_out_Y       , B1, and0_out          );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__A21OI_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__A21OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a21oi: 2-input AND into first input of 2-input NOR.
 *
 *        Y = !((A1 & A2) | B1)
 *
 * Verilog wrapper for a21oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__a21oi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__a21oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__A21OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22o: 2-input AND into both inputs of 2-input OR.
 *
 *       X = ((A1 & A2) | (B1 & B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a22o: 2-input AND into both inputs of 2-input OR.
 *
 *       X = ((A1 & A2) | (B1 & B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__a22o (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out         ;
    wire and1_out         ;
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    and                                 and0        (and0_out         , B1, B2               );
    and                                 and1        (and1_out         , A1, A2               );
    or                                  or0         (or0_out_X        , and1_out, and0_out   );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__A22O_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__A22O_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22o: 2-input AND into both inputs of 2-input OR.
 *
 *       X = ((A1 & A2) | (B1 & B2))
 *
 * Verilog wrapper for a22o with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__a22o_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__a22o base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__A22O_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22oi: 2-input AND into both inputs of 2-input NOR.
 *
 *        Y = !((A1 & A2) | (B1 & B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * a22oi: 2-input AND into both inputs of 2-input NOR.
 *
 *        Y = !((A1 & A2) | (B1 & B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__a22oi (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out        ;
    wire nand1_out        ;
    wire and0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    nand                                nand0       (nand0_out        , A2, A1                );
    nand                                nand1       (nand1_out        , B2, B1                );
    and                                 and0        (and0_out_Y       , nand0_out, nand1_out  );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, and0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__A22OI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__A22OI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * a22oi: 2-input AND into both inputs of 2-input NOR.
 *
 *        Y = !((A1 & A2) | (B1 & B2))
 *
 * Verilog wrapper for a22oi with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__a22oi_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__a22oi base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__A22OI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2: 2-input AND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and2: 2-input AND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__and2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    and                                 and0        (and0_out_X       , A, B                  );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__AND2_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__AND2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and2: 2-input AND.
 *
 * Verilog wrapper for and2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__and2_1 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__and2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__AND2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3: 3-input AND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * and3: 3-input AND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__and3 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    and                                 and0        (and0_out_X       , C, A, B               );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__AND3_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__AND3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * and3: 3-input AND.
 *
 * Verilog wrapper for and3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__and3_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__and3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__AND3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * buf: Buffer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__buf (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    buf                                 buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                 buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__BUF_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__BUF_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__buf_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__BUF_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__buf_2 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__BUF_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__buf_4 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__BUF_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__buf_8 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__BUF_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__buf_16 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__BUF_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * buf: Buffer.
 *
 * Verilog wrapper for buf with size of 32 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__buf_32 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__buf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__BUF_32_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * conb: Constant value, low, high outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * conb: Constant value, low, high outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__conb (
    HI  ,
    LO  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output HI  ;
    output LO  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire pullup0_out_HI  ;
    wire pulldown0_out_LO;

    //                                 Name         Output            Other arguments
    pullup                             pullup0     (pullup0_out_HI  );
    sky130_fd_sc_hvl__udp_pwrgood_pp$P pwrgood_pp0 (HI              , pullup0_out_HI, VPWR  );
    pulldown                           pulldown0   (pulldown0_out_LO);
    sky130_fd_sc_hvl__udp_pwrgood_pp$G pwrgood_pp1 (LO              , pulldown0_out_LO, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__CONB_FUNCTIONAL_PP_V



































































 // FUNCTIONAL

















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__CONB_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * conb: Constant value, low, high outputs.
 *
 * Verilog wrapper for conb with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__conb_1 (
    HI  ,
    LO  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output HI  ;
    output LO  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__conb base (
        .HI(HI),
        .LO(LO),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__CONB_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hvl__decap (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DECAP_FUNCTIONAL_PP_V



















































 // FUNCTIONAL



























































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DECAP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog wrapper for decap with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__decap_4 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hvl__decap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DECAP_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * decap: Decoupling capacitance filler.
 *
 * Verilog wrapper for decap with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__decap_8 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hvl__decap base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DECAP_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrbp: Delay flop, inverted reset, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfrbp: Delay flop, inverted reset, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dfrbp (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q      ;
    wire RESET      ;
    wire buf0_out_Q ;
    wire not1_out_qn;

    //                                   Delay       Name         Output       Other arguments
    not                                              not0        (RESET      , RESET_B                    );
    sky130_fd_sc_hvl__udp_dff$PR_pp$PG$N #1 dff0        (buf_Q      , D, CLK, RESET, , VPWR, VGND);
    buf                                              buf0        (buf0_out_Q , buf_Q                      );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp0 (Q          , buf0_out_Q, VPWR, VGND     );
    not                                              not1        (not1_out_qn, buf_Q                      );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp1 (Q_N        , not1_out_qn, VPWR, VGND    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DFRBP_FUNCTIONAL_PP_V



















































































 // FUNCTIONAL



















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFRBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrbp: Delay flop, inverted reset, complementary outputs.
 *
 * Verilog wrapper for dfrbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dfrbp_1 (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hvl__dfrbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFRBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrtp: Delay flop, inverted reset, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfrtp: Delay flop, inverted reset, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dfrtp (
    Q      ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q     ;
    wire RESET     ;
    wire buf0_out_Q;

    //                                   Delay       Name         Output      Other arguments
    not                                              not0        (RESET     , RESET_B                    );
    sky130_fd_sc_hvl__udp_dff$PR_pp$PG$N #1 dff0        (buf_Q     , D, CLK, RESET, , VPWR, VGND);
    buf                                              buf0        (buf0_out_Q, buf_Q                      );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DFRTP_FUNCTIONAL_PP_V














































































 // FUNCTIONAL













































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFRTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfrtp: Delay flop, inverted reset, single output.
 *
 * Verilog wrapper for dfrtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dfrtp_1 (
    Q      ,
    CLK    ,
    D      ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK    ;
    input  D      ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hvl__dfrtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFRTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfsbp: Delay flop, inverted set, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfsbp: Delay flop, inverted set, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dfsbp (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf_Q      ;
    wire SET        ;
    wire buf0_out_Q ;
    wire not1_out_qn;

    //                                   Delay       Name         Output       Other arguments
    not                                              not0        (SET        , SET_B                    );
    sky130_fd_sc_hvl__udp_dff$PS_pp$PG$N #1 dff0        (buf_Q      , D, CLK, SET, , VPWR, VGND);
    buf                                              buf0        (buf0_out_Q , buf_Q                    );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp0 (Q          , buf0_out_Q, VPWR, VGND   );
    not                                              not1        (not1_out_qn, buf_Q                    );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp1 (Q_N        , not1_out_qn, VPWR, VGND  );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DFSBP_FUNCTIONAL_PP_V



















































































 // FUNCTIONAL



















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFSBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfsbp: Delay flop, inverted set, complementary outputs.
 *
 * Verilog wrapper for dfsbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dfsbp_1 (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hvl__dfsbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFSBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfstp: Delay flop, inverted set, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfstp: Delay flop, inverted set, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dfstp (
    Q    ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf_Q     ;
    wire SET       ;
    wire buf0_out_Q;

    //                                   Delay       Name         Output      Other arguments
    not                                              not0        (SET       , SET_B                    );
    sky130_fd_sc_hvl__udp_dff$PS_pp$PG$N #1 dff0        (buf_Q     , D, CLK, SET, , VPWR, VGND);
    buf                                              buf0        (buf0_out_Q, buf_Q                    );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND   );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DFSTP_FUNCTIONAL_PP_V














































































 // FUNCTIONAL













































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFSTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfstp: Delay flop, inverted set, single output.
 *
 * Verilog wrapper for dfstp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dfstp_1 (
    Q    ,
    CLK  ,
    D    ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hvl__dfstp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFSTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxbp: Delay flop, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfxbp: Delay flop, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dfxbp (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q      ;
    wire buf0_out_Q ;
    wire not0_out_qn;

    //                                  Delay       Name         Output       Other arguments
    sky130_fd_sc_hvl__udp_dff$P_pp$PG$N #1 dff0        (buf_Q      , D, CLK, , VPWR, VGND   );
    buf                                             buf0        (buf0_out_Q , buf_Q                  );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG             pwrgood_pp0 (Q          , buf0_out_Q, VPWR, VGND );
    not                                             not0        (not0_out_qn, buf_Q                  );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG             pwrgood_pp1 (Q_N        , not0_out_qn, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DFXBP_FUNCTIONAL_PP_V












































































 // FUNCTIONAL








































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFXBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxbp: Delay flop, complementary outputs.
 *
 * Verilog wrapper for dfxbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dfxbp_1 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__dfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFXBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxtp: Delay flop, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dfxtp: Delay flop, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dfxtp (
    Q   ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q     ;
    wire buf0_out_Q;

    //                                  Delay       Name         Output      Other arguments
    sky130_fd_sc_hvl__udp_dff$P_pp$PG$N #1 dff0        (buf_Q     , D, CLK, , VPWR, VGND  );
    buf                                             buf0        (buf0_out_Q, buf_Q                 );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG             pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DFXTP_FUNCTIONAL_PP_V







































































 // FUNCTIONAL


































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dfxtp: Delay flop, single output.
 *
 * Verilog wrapper for dfxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dfxtp_1 (
    Q   ,
    CLK ,
    D   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__dfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DFXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * diode: Antenna tie-down diode.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * diode: Antenna tie-down diode.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hvl__diode (
    DIODE,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    input DIODE;
    input VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DIODE_FUNCTIONAL_PP_V





















































 // FUNCTIONAL





































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DIODE_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * diode: Antenna tie-down diode.
 *
 * Verilog wrapper for diode with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__diode_2 (
    DIODE,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    input DIODE;
    input VPWR ;
    input VGND ;
    input VPB  ;
    input VNB  ;
    sky130_fd_sc_hvl__diode base (
        .DIODE(DIODE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/
























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DIODE_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlclkp: Clock gate.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlclkp: Clock gate.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dlclkp (
    GCLK,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output GCLK;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire m0    ;
    wire clkn  ;
    wire GCLK_b;

    //                                     Name         Output  Other arguments
    not                                    not0        (clkn  , CLK                     );
    sky130_fd_sc_hvl__udp_dlatch$P_pp$PG$N dlatch0     (m0    , GATE, clkn, , VPWR, VGND);
    and                                    and0        (GCLK_b, m0, CLK                 );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG    pwrgood_pp0 (GCLK  , GCLK_b, VPWR, VGND      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DLCLKP_FUNCTIONAL_PP_V











































































 // FUNCTIONAL










































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DLCLKP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlclkp: Clock gate.
 *
 * Verilog wrapper for dlclkp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dlclkp_1 (
    GCLK,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output GCLK;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__dlclkp base (
        .GCLK(GCLK),
        .GATE(GATE),
        .CLK(CLK),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DLCLKP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtp: Delay latch, inverted reset, non-inverted enable,
 *        single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlrtp: Delay latch, inverted reset, non-inverted enable,
 *        single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dlrtp (
    Q      ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire RESET     ;
    wire buf_Q     ;
    wire buf0_out_Q;

    //                                      Delay       Name         Output      Other arguments
    not                                                 not0        (RESET     , RESET_B                     );
    sky130_fd_sc_hvl__udp_dlatch$PR_pp$PG$N #1 dlatch0     (buf_Q     , D, GATE, RESET, , VPWR, VGND);
    buf                                                 buf0        (buf0_out_Q, buf_Q                       );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG                 pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DLRTP_FUNCTIONAL_PP_V
















































































 // FUNCTIONAL
















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DLRTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlrtp: Delay latch, inverted reset, non-inverted enable,
 *        single output.
 *
 * Verilog wrapper for dlrtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dlrtp_1 (
    Q      ,
    RESET_B,
    D      ,
    GATE   ,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  RESET_B;
    input  D      ;
    input  GATE   ;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hvl__dlrtp base (
        .Q(Q),
        .RESET_B(RESET_B),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DLRTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxtp: Delay latch, non-inverted enable, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * dlxtp: Delay latch, non-inverted enable, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__dlxtp (
    Q   ,
    D   ,
    GATE,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  D   ;
    input  GATE;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q     ;
    wire buf0_out_Q;

    //                                     Delay       Name         Output      Other arguments
    sky130_fd_sc_hvl__udp_dlatch$P_pp$PG$N #1 dlatch0     (buf_Q     , D, GATE, , VPWR, VGND );
    buf                                                buf0        (buf0_out_Q, buf_Q                 );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG                pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__DLXTP_FUNCTIONAL_PP_V







































































 // FUNCTIONAL


































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DLXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * dlxtp: Delay latch, non-inverted enable, single output.
 *
 * Verilog wrapper for dlxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__dlxtp_1 (
    Q   ,
    D   ,
    GATE,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  D   ;
    input  GATE;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__dlxtp base (
        .Q(Q),
        .D(D),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__DLXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__einvn (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire pwrgood_pp0_out_A  ;
    wire pwrgood_pp1_out_teb;

    //                                  Name         Output               Other arguments
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A  , A, VPWR, VGND                         );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_teb, TE_B, VPWR, VGND                      );
    notif0                              notif00     (Z                  , pwrgood_pp0_out_A, pwrgood_pp1_out_teb);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__EINVN_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__EINVN_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvn: Tri-state inverter, negative enable.
 *
 * Verilog wrapper for einvn with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__einvn_1 (
    Z   ,
    A   ,
    TE_B,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE_B;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__einvn base (
        .Z(Z),
        .A(A),
        .TE_B(TE_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__EINVN_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__einvp (
    Z   ,
    A   ,
    TE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Z   ;
    input  A   ;
    input  TE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire pwrgood_pp0_out_A ;
    wire pwrgood_pp1_out_TE;

    //                                  Name         Output              Other arguments
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A , A, VPWR, VGND                        );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp1 (pwrgood_pp1_out_TE, TE, VPWR, VGND                       );
    notif1                              notif10     (Z                 , pwrgood_pp0_out_A, pwrgood_pp1_out_TE);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__EINVP_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__EINVP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * einvp: Tri-state inverter, positive enable.
 *
 * Verilog wrapper for einvp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__einvp_1 (
    Z   ,
    A   ,
    TE  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Z   ;
    input  A   ;
    input  TE  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__einvp base (
        .Z(Z),
        .A(A),
        .TE(TE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__EINVP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * fill: Fill cell.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_hvl__fill (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
     // No contents.
endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__FILL_FUNCTIONAL_PP_V



















































 // FUNCTIONAL

































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__FILL_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__fill_1 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hvl__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__FILL_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__fill_2 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hvl__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__FILL_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__fill_4 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hvl__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__FILL_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * fill: Fill cell.
 *
 * Verilog wrapper for fill with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__fill_8 (
    VPWR,
    VGND,
    VPB ,
    VNB
);

    input VPWR;
    input VGND;
    input VPB ;
    input VNB ;
    sky130_fd_sc_hvl__fill base (
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

















 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__FILL_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * inv: Inverter.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__inv (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire not0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    not                                 not0        (not0_out_Y       , A                     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, not0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__INV_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__INV_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__inv_1 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__INV_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 2 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__inv_2 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__INV_2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 4 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__inv_4 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__INV_4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__inv_8 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__INV_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * inv: Inverter.
 *
 * Verilog wrapper for inv with size of 16 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__inv_16 (
    Y   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__inv base (
        .Y(Y),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__INV_16_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbufhv2hv_hl: Level shifting buffer, High Voltage to High Voltage,
 *                Higher Voltage to Lower Voltage.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lsbufhv2hv_hl: Level shifting buffer, High Voltage to High Voltage,
 *                Higher Voltage to Lower Voltage.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__lsbufhv2hv_hl (
    X       ,
    A       ,
    VPWR    ,
    VGND    ,
    LOWHVPWR,
    VPB     ,
    VNB
);

    // Module ports
    output X       ;
    input  A       ;
    input  VPWR    ;
    input  VGND    ;
    input  LOWHVPWR;
    input  VPB     ;
    input  VNB     ;

    // Local signals
    wire pwrgood_pp0_out_A;
    wire buf0_out_X       ;

    //                                  Name         Output             Other arguments
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A, A, VPWR, VGND             );
    buf                                 buf0        (buf0_out_X       , pwrgood_pp0_out_A         );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp1 (X                , buf0_out_X, LOWHVPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2HV_HL_FUNCTIONAL_PP_V





































































 // FUNCTIONAL


















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2HV_HL_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbufhv2hv_hl: Level shifting buffer, High Voltage to High Voltage,
 *                Higher Voltage to Lower Voltage.
 *
 * Verilog wrapper for lsbufhv2hv_hl with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__lsbufhv2hv_hl_1 (
    X       ,
    A       ,
    VPWR    ,
    VGND    ,
    LOWHVPWR,
    VPB     ,
    VNB
);

    output X       ;
    input  A       ;
    input  VPWR    ;
    input  VGND    ;
    input  LOWHVPWR;
    input  VPB     ;
    input  VNB     ;
    sky130_fd_sc_hvl__lsbufhv2hv_hl base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .LOWHVPWR(LOWHVPWR),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbufhv2hv_lh: Level shifting buffer, High Voltage to High Voltage,
 *                Lower Voltage to Higher Voltage.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lsbufhv2hv_lh: Level shifting buffer, High Voltage to High Voltage,
 *                Lower Voltage to Higher Voltage.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__lsbufhv2hv_lh (
    X       ,
    A       ,
    VPWR    ,
    VGND    ,
    LOWHVPWR,
    VPB     ,
    VNB
);

    // Module ports
    output X       ;
    input  A       ;
    input  VPWR    ;
    input  VGND    ;
    input  LOWHVPWR;
    input  VPB     ;
    input  VNB     ;

    // Local signals
    wire pwrgood_pp0_out_A;
    wire buf0_out_X       ;

    //                                  Name         Output             Other arguments
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A, A, LOWHVPWR, VGND     );
    buf                                 buf0        (buf0_out_X       , pwrgood_pp0_out_A     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp1 (X                , buf0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2HV_LH_FUNCTIONAL_PP_V





































































 // FUNCTIONAL


















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2HV_LH_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbufhv2hv_lh: Level shifting buffer, High Voltage to High Voltage,
 *                Lower Voltage to Higher Voltage.
 *
 * Verilog wrapper for lsbufhv2hv_lh with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__lsbufhv2hv_lh_1 (
    X       ,
    A       ,
    VPWR    ,
    VGND    ,
    LOWHVPWR,
    VPB     ,
    VNB
);

    output X       ;
    input  A       ;
    input  VPWR    ;
    input  VGND    ;
    input  LOWHVPWR;
    input  VPB     ;
    input  VNB     ;
    sky130_fd_sc_hvl__lsbufhv2hv_lh base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .LOWHVPWR(LOWHVPWR),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbufhv2lv: Level-shift buffer, low voltage-to-low voltage.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lsbufhv2lv: Level-shift buffer, low voltage-to-low voltage.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__lsbufhv2lv (
    X    ,
    A    ,
    VPWR ,
    VGND ,
    LVPWR,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  LVPWR;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire pwrgood_pp0_out_A;
    wire buf0_out_X       ;

    //                                  Name         Output             Other arguments
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A, A, VPWR, VGND          );
    buf                                 buf0        (buf0_out_X       , pwrgood_pp0_out_A      );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp1 (X                , buf0_out_X, LVPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2LV_FUNCTIONAL_PP_V




































































 // FUNCTIONAL
















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2LV_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbufhv2lv: Level-shift buffer, low voltage-to-low voltage.
 *
 * Verilog wrapper for lsbufhv2lv with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__lsbufhv2lv_1 (
    X    ,
    A    ,
    VPWR ,
    VGND ,
    LVPWR,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  LVPWR;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hvl__lsbufhv2lv base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .LVPWR(LVPWR),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2LV_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbufhv2lv_simple: Level shifting buffer, High Voltage to Low
 *                    Voltage, simple (hv devices in inverters on lv
 *                    power rail).
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lsbufhv2lv_simple: Level shifting buffer, High Voltage to Low
 *                    Voltage, simple (hv devices in inverters on lv
 *                    power rail).
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__lsbufhv2lv_simple (
    X    ,
    A    ,
    VPWR ,
    VGND ,
    LVPWR,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  LVPWR;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire pwrgood_pp0_out_A;
    wire buf0_out_X       ;

    //                                  Name         Output             Other arguments
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A, A, VPWR, VGND          );
    buf                                 buf0        (buf0_out_X       , pwrgood_pp0_out_A      );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp1 (X                , buf0_out_X, LVPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_FUNCTIONAL_PP_V






































































 // FUNCTIONAL




















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbufhv2lv_simple: Level shifting buffer, High Voltage to Low
 *                    Voltage, simple (hv devices in inverters on lv
 *                    power rail).
 *
 * Verilog wrapper for lsbufhv2lv_simple with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__lsbufhv2lv_simple_1 (
    X    ,
    A    ,
    VPWR ,
    VGND ,
    LVPWR,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  LVPWR;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hvl__lsbufhv2lv_simple base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .LVPWR(LVPWR),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbuflv2hv: Level-shift buffer, low voltage-to-high voltage,
 *             isolated well on input buffer, double height cell.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lsbuflv2hv: Level-shift buffer, low voltage-to-high voltage,
 *             isolated well on input buffer, double height cell.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__lsbuflv2hv (
    X    ,
    A    ,
    VPWR ,
    VGND ,
    LVPWR,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  LVPWR;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire pwrgood_pp0_out_A;
    wire buf0_out_X       ;

    //                                  Name         Output             Other arguments
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A, A, LVPWR, VGND        );
    buf                                 buf0        (buf0_out_X       , pwrgood_pp0_out_A     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp1 (X                , buf0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_FUNCTIONAL_PP_V





































































 // FUNCTIONAL


















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbuflv2hv: Level-shift buffer, low voltage-to-high voltage,
 *             isolated well on input buffer, double height cell.
 *
 * Verilog wrapper for lsbuflv2hv with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__lsbuflv2hv_1 (
    X    ,
    A    ,
    VPWR ,
    VGND ,
    LVPWR,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  LVPWR;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hvl__lsbuflv2hv base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .LVPWR(LVPWR),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbuflv2hv_clkiso_hlkg: Level-shift clock buffer, low voltage to
 *                         high voltage, isolated well
 *                         on input buffer, inverting sleep
 *                         mode input.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lsbuflv2hv_clkiso_hlkg: Level-shift clock buffer, low voltage to
 *                         high voltage, isolated well
 *                         on input buffer, inverting sleep
 *                         mode input.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg (
    X      ,
    A      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    LVPWR  ,
    VPB    ,
    VNB
);

    // Module ports
    output X      ;
    input  A      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  LVPWR  ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire SLEEP               ;
    wire and0_out_X          ;
    wire isolatchhv_pp0_out_X;

    //                                        Name            Output                Other arguments
    not                                       not0           (SLEEP               , SLEEP_B                             );
    and                                       and0           (and0_out_X          , SLEEP_B, A                          );
    sky130_fd_sc_hvl__udp_isolatchhv_pp$PLG$S isolatchhv_pp0 (isolatchhv_pp0_out_X, and0_out_X, VPWR, LVPWR, VGND, SLEEP);
    buf                                       buf0           (X                   , isolatchhv_pp0_out_X                );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_FUNCTIONAL_PP_V











































































 // FUNCTIONAL






































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbuflv2hv_clkiso_hlkg: Level-shift clock buffer, low voltage to
 *                         high voltage, isolated well
 *                         on input buffer, inverting sleep
 *                         mode input.
 *
 * Verilog wrapper for lsbuflv2hv_clkiso_hlkg with size of 3 units
 * (invalid?).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3 (
    X      ,
    A      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    LVPWR  ,
    VPB    ,
    VNB
);

    output X      ;
    input  A      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  LVPWR  ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg base (
        .X(X),
        .A(A),
        .SLEEP_B(SLEEP_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .LVPWR(LVPWR),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbuflv2hv_isosrchvaon: Level shift buffer, low voltage to high
 *                         voltage, isolated well on input buffer,
 *                         inverting sleep mode input, zero power
 *                         sleep mode.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lsbuflv2hv_isosrchvaon: Level shift buffer, low voltage to high
 *                         voltage, isolated well on input buffer,
 *                         inverting sleep mode input, zero power
 *                         sleep mode.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon (
    X      ,
    A      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    LVPWR  ,
    VPB    ,
    VNB
);

    // Module ports
    output X      ;
    input  A      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  LVPWR  ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire SLEEP               ;
    wire and0_out_X          ;
    wire isolatchhv_pp0_out_X;

    //                                        Name            Output                Other arguments
    not                                       not0           (SLEEP               , SLEEP_B                             );
    and                                       and0           (and0_out_X          , SLEEP_B, A                          );
    sky130_fd_sc_hvl__udp_isolatchhv_pp$PLG$S isolatchhv_pp0 (isolatchhv_pp0_out_X, and0_out_X, VPWR, LVPWR, VGND, SLEEP);
    buf                                       buf0           (X                   , isolatchhv_pp0_out_X                );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_FUNCTIONAL_PP_V











































































 // FUNCTIONAL






































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbuflv2hv_isosrchvaon: Level shift buffer, low voltage to high
 *                         voltage, isolated well on input buffer,
 *                         inverting sleep mode input, zero power
 *                         sleep mode.
 *
 * Verilog wrapper for lsbuflv2hv_isosrchvaon with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1 (
    X      ,
    A      ,
    SLEEP_B,
    VPWR   ,
    VGND   ,
    LVPWR  ,
    VPB    ,
    VNB
);

    output X      ;
    input  A      ;
    input  SLEEP_B;
    input  VPWR   ;
    input  VGND   ;
    input  LVPWR  ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon base (
        .X(X),
        .A(A),
        .SLEEP_B(SLEEP_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .LVPWR(LVPWR),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbuflv2hv_symmetric: Level shifting buffer, Low Voltage to High
 *                       Voltage, Symmetrical.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * lsbuflv2hv_symmetric: Level shifting buffer, Low Voltage to High
 *                       Voltage, Symmetrical.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__lsbuflv2hv_symmetric (
    X    ,
    A    ,
    VPWR ,
    VGND ,
    LVPWR,
    VPB  ,
    VNB
);

    // Module ports
    output X    ;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  LVPWR;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire pwrgood_pp0_out_A;
    wire buf0_out_X       ;

    //                                  Name         Output             Other arguments
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_A, A, LVPWR, VGND        );
    buf                                 buf0        (buf0_out_X       , pwrgood_pp0_out_A     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp1 (X                , buf0_out_X, VPWR, VGND);

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_FUNCTIONAL_PP_V





































































 // FUNCTIONAL


















































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * lsbuflv2hv_symmetric: Level shifting buffer, Low Voltage to High
 *                       Voltage, Symmetrical.
 *
 * Verilog wrapper for lsbuflv2hv_symmetric with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1 (
    X    ,
    A    ,
    VPWR ,
    VGND ,
    LVPWR,
    VPB  ,
    VNB
);

    output X    ;
    input  A    ;
    input  VPWR ;
    input  VGND ;
    input  LVPWR;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hvl__lsbuflv2hv_symmetric base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .LVPWR(LVPWR),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2: 2-input multiplexer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * mux2: 2-input multiplexer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__mux2 (
    X   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire mux_2to10_out_X  ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    sky130_fd_sc_hvl__udp_mux_2to1      mux_2to10   (mux_2to10_out_X  , A0, A1, S                  );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, mux_2to10_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__MUX2_FUNCTIONAL_PP_V






































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__MUX2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux2: 2-input multiplexer.
 *
 * Verilog wrapper for mux2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__mux2_1 (
    X   ,
    A0  ,
    A1  ,
    S   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  S   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__mux2 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .S(S),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__MUX2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux4: 4-input multiplexer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * mux4: 4-input multiplexer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__mux4 (
    X   ,
    A0  ,
    A1  ,
    A2  ,
    A3  ,
    S0  ,
    S1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A0  ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  S0  ;
    input  S1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire mux_4to20_out_X  ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    sky130_fd_sc_hvl__udp_mux_4to2      mux_4to20   (mux_4to20_out_X  , A0, A1, A2, A3, S0, S1     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, mux_4to20_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__MUX4_FUNCTIONAL_PP_V












































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__MUX4_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * mux4: 4-input multiplexer.
 *
 * Verilog wrapper for mux4 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__mux4_1 (
    X   ,
    A0  ,
    A1  ,
    A2  ,
    A3  ,
    S0  ,
    S1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A0  ;
    input  A1  ;
    input  A2  ;
    input  A3  ;
    input  S0  ;
    input  S1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__mux4 base (
        .X(X),
        .A0(A0),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .S0(S0),
        .S1(S1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__MUX4_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2: 2-input NAND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand2: 2-input NAND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__nand2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    nand                                nand0       (nand0_out_Y      , B, A                   );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__NAND2_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__NAND2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand2: 2-input NAND.
 *
 * Verilog wrapper for nand2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__nand2_1 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__nand2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__NAND2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3: 3-input NAND.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nand3: 3-input NAND.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__nand3 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    nand                                nand0       (nand0_out_Y      , B, A, C                );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__NAND3_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__NAND3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nand3: 3-input NAND.
 *
 * Verilog wrapper for nand3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__nand3_1 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__nand3 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__NAND3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2: 2-input NOR.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor2: 2-input NOR.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__nor2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    nor                                 nor0        (nor0_out_Y       , A, B                  );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__NOR2_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__NOR2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor2: 2-input NOR.
 *
 * Verilog wrapper for nor2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__nor2_1 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__nor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__NOR2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3: 3-input NOR.
 *
 *       Y = !(A | B | C | !D)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * nor3: 3-input NOR.
 *
 *       Y = !(A | B | C | !D)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__nor3 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out_Y       ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    nor                                 nor0        (nor0_out_Y       , C, A, B               );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nor0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__NOR3_FUNCTIONAL_PP_V








































































 // FUNCTIONAL



































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__NOR3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * nor3: 3-input NOR.
 *
 *       Y = !(A | B | C | !D)
 *
 * Verilog wrapper for nor3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__nor3_1 (
    Y   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__nor3 base (
        .Y(Y),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__NOR3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21a: 2-input OR into first input of 2-input AND.
 *
 *       X = ((A1 | A2) & B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o21a: 2-input OR into first input of 2-input AND.
 *
 *       X = ((A1 | A2) & B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__o21a (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    or                                  or0         (or0_out          , A2, A1                );
    and                                 and0        (and0_out_X       , or0_out, B1           );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__O21A_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__O21A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21a: 2-input OR into first input of 2-input AND.
 *
 *       X = ((A1 | A2) & B1)
 *
 * Verilog wrapper for o21a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__o21a_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__o21a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__O21A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__o21ai (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire nand0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    or                                  or0         (or0_out          , A2, A1                 );
    nand                                nand0       (nand0_out_Y      , B1, or0_out            );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, nand0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__O21AI_FUNCTIONAL_PP_V










































































 // FUNCTIONAL







































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__O21AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o21ai: 2-input OR into first input of 2-input NAND.
 *
 *        Y = !((A1 | A2) & B1)
 *
 * Verilog wrapper for o21ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__o21ai_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__o21ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__O21AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22a: 2-input OR into both inputs of 2-input AND.
 *
 *       X = ((A1 | A2) & (B1 | B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o22a: 2-input OR into both inputs of 2-input AND.
 *
 *       X = ((A1 | A2) & (B1 | B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__o22a (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out          ;
    wire or1_out          ;
    wire and0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    or                                  or0         (or0_out          , A2, A1                );
    or                                  or1         (or1_out          , B2, B1                );
    and                                 and0        (and0_out_X       , or0_out, or1_out      );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, and0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__O22A_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__O22A_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22a: 2-input OR into both inputs of 2-input AND.
 *
 *       X = ((A1 | A2) & (B1 | B2))
 *
 * Verilog wrapper for o22a with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__o22a_1 (
    X   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__o22a base (
        .X(X),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__O22A_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22ai: 2-input OR into both inputs of 2-input NAND.
 *
 *        Y = !((A1 | A2) & (B1 | B2))
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * o22ai: 2-input OR into both inputs of 2-input NAND.
 *
 *        Y = !((A1 | A2) & (B1 | B2))
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__o22ai (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire nor0_out         ;
    wire nor1_out         ;
    wire or0_out_Y        ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    nor                                 nor0        (nor0_out         , B1, B2               );
    nor                                 nor1        (nor1_out         , A1, A2               );
    or                                  or0         (or0_out_Y        , nor1_out, nor0_out   );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, or0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__O22AI_FUNCTIONAL_PP_V














































































 // FUNCTIONAL















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__O22AI_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * o22ai: 2-input OR into both inputs of 2-input NAND.
 *
 *        Y = !((A1 | A2) & (B1 | B2))
 *
 * Verilog wrapper for o22ai with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__o22ai_1 (
    Y   ,
    A1  ,
    A2  ,
    B1  ,
    B2  ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A1  ;
    input  A2  ;
    input  B1  ;
    input  B2  ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__o22ai base (
        .Y(Y),
        .A1(A1),
        .A2(A2),
        .B1(B1),
        .B2(B2),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__O22AI_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2: 2-input OR.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or2: 2-input OR.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__or2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    or                                  or0         (or0_out_X        , B, A                 );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__OR2_FUNCTIONAL_PP_V




































































 // FUNCTIONAL



























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__OR2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or2: 2-input OR.
 *
 * Verilog wrapper for or2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__or2_1 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__or2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__OR2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3: 3-input OR.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * or3: 3-input OR.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__or3 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire or0_out_X        ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    or                                  or0         (or0_out_X        , B, A, C              );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, or0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__OR3_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__OR3_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * or3: 3-input OR.
 *
 * Verilog wrapper for or3 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__or3_1 (
    X   ,
    A   ,
    B   ,
    C   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__or3 base (
        .X(X),
        .A(A),
        .B(B),
        .C(C),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__OR3_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * probe_p: Virtual voltage probe point.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * probe_p: Virtual voltage probe point.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__probe_p (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    buf                                 buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                 buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__PROBE_P_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__PROBE_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * probe_p: Virtual voltage probe point.
 *
 * Verilog wrapper for probe_p with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__probe_p_8 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__probe_p base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__PROBE_P_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * probec_p: Virtual current probe point.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * probec_p: Virtual current probe point.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__probec_p (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    buf                                 buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                 buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__PROBEC_P_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__PROBEC_P_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * probec_p: Virtual current probe point.
 *
 * Verilog wrapper for probec_p with size of 8 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__probec_p_8 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__probec_p base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__PROBEC_P_8_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * schmittbuf: Schmitt Trigger Buffer.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * schmittbuf: Schmitt Trigger Buffer.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__schmittbuf (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    buf                                 buf0        (buf0_out_X       , A                     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, buf0_out_X, VPWR, VGND);
    buf                                 buf1        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SCHMITTBUF_FUNCTIONAL_PP_V


































































 // FUNCTIONAL























































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SCHMITTBUF_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * schmittbuf: Schmitt Trigger Buffer.
 *
 * Verilog wrapper for schmittbuf with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__schmittbuf_1 (
    X   ,
    A   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__schmittbuf base (
        .X(X),
        .A(A),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/



























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SCHMITTBUF_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrbp: Scan delay flop, inverted reset, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfrbp: Scan delay flop, inverted reset, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__sdfrbp (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q      ;
    wire RESET      ;
    wire mux_out    ;
    wire buf0_out_Q ;
    wire not1_out_qn;

    //                                   Delay       Name         Output       Other arguments
    not                                              not0        (RESET      , RESET_B                          );
    sky130_fd_sc_hvl__udp_mux_2to1                   mux_2to10   (mux_out    , D, SCD, SCE                      );
    sky130_fd_sc_hvl__udp_dff$PR_pp$PG$N #1 dff0        (buf_Q      , mux_out, CLK, RESET, , VPWR, VGND);
    buf                                              buf0        (buf0_out_Q , buf_Q                            );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp0 (Q          , buf0_out_Q, VPWR, VGND           );
    not                                              not1        (not1_out_qn, buf_Q                            );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp1 (Q_N        , not1_out_qn, VPWR, VGND          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFRBP_FUNCTIONAL_PP_V


































































































 // FUNCTIONAL









































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFRBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrbp: Scan delay flop, inverted reset, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog wrapper for sdfrbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__sdfrbp_1 (
    Q      ,
    Q_N    ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    output Q_N    ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hvl__sdfrbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFRBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrtp: Scan delay flop, inverted reset, non-inverted clock,
 *         single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfrtp: Scan delay flop, inverted reset, non-inverted clock,
 *         single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__sdfrtp (
    Q      ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    // Module ports
    output Q      ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;

    // Local signals
    wire buf_Q     ;
    wire RESET     ;
    wire mux_out   ;
    wire buf0_out_Q;

    //                                   Delay       Name         Output      Other arguments
    not                                              not0        (RESET     , RESET_B                          );
    sky130_fd_sc_hvl__udp_mux_2to1                   mux_2to10   (mux_out   , D, SCD, SCE                      );
    sky130_fd_sc_hvl__udp_dff$PR_pp$PG$N #1 dff0        (buf_Q     , mux_out, CLK, RESET, , VPWR, VGND);
    buf                                              buf0        (buf0_out_Q, buf_Q                            );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND           );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFRTP_FUNCTIONAL_PP_V





























































































 // FUNCTIONAL



































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFRTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfrtp: Scan delay flop, inverted reset, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfrtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__sdfrtp_1 (
    Q      ,
    CLK    ,
    D      ,
    SCD    ,
    SCE    ,
    RESET_B,
    VPWR   ,
    VGND   ,
    VPB    ,
    VNB
);

    output Q      ;
    input  CLK    ;
    input  D      ;
    input  SCD    ;
    input  SCE    ;
    input  RESET_B;
    input  VPWR   ;
    input  VGND   ;
    input  VPB    ;
    input  VNB    ;
    sky130_fd_sc_hvl__sdfrtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .RESET_B(RESET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFRTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfsbp: Scan delay flop, inverted set, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfsbp: Scan delay flop, inverted set, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__sdfsbp (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf_Q      ;
    wire SET        ;
    wire mux_out    ;
    wire buf0_out_Q ;
    wire not1_out_qn;

    //                                   Delay       Name         Output       Other arguments
    not                                              not0        (SET        , SET_B                          );
    sky130_fd_sc_hvl__udp_mux_2to1                   mux_2to10   (mux_out    , D, SCD, SCE                    );
    sky130_fd_sc_hvl__udp_dff$PS_pp$PG$N #1 dff0        (buf_Q      , mux_out, CLK, SET, , VPWR, VGND);
    buf                                              buf0        (buf0_out_Q , buf_Q                          );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp0 (Q          , buf0_out_Q, VPWR, VGND         );
    not                                              not1        (not1_out_qn, buf_Q                          );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp1 (Q_N        , not1_out_qn, VPWR, VGND        );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFSBP_FUNCTIONAL_PP_V


































































































 // FUNCTIONAL









































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFSBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfsbp: Scan delay flop, inverted set, non-inverted clock,
 *         complementary outputs.
 *
 * Verilog wrapper for sdfsbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__sdfsbp_1 (
    Q    ,
    Q_N  ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    output Q_N  ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hvl__sdfsbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/










































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFSBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfstp: Scan delay flop, inverted set, non-inverted clock,
 *         single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfstp: Scan delay flop, inverted set, non-inverted clock,
 *         single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__sdfstp (
    Q    ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    // Module ports
    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;

    // Local signals
    wire buf_Q     ;
    wire SET       ;
    wire mux_out   ;
    wire buf0_out_Q;

    //                                   Delay       Name         Output      Other arguments
    not                                              not0        (SET       , SET_B                          );
    sky130_fd_sc_hvl__udp_mux_2to1                   mux_2to10   (mux_out   , D, SCD, SCE                    );
    sky130_fd_sc_hvl__udp_dff$PS_pp$PG$N #1 dff0        (buf_Q     , mux_out, CLK, SET, , VPWR, VGND);
    buf                                              buf0        (buf0_out_Q, buf_Q                          );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG              pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND         );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFSTP_FUNCTIONAL_PP_V





























































































 // FUNCTIONAL



































































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFSTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfstp: Scan delay flop, inverted set, non-inverted clock,
 *         single output.
 *
 * Verilog wrapper for sdfstp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__sdfstp_1 (
    Q    ,
    CLK  ,
    D    ,
    SCD  ,
    SCE  ,
    SET_B,
    VPWR ,
    VGND ,
    VPB  ,
    VNB
);

    output Q    ;
    input  CLK  ;
    input  D    ;
    input  SCD  ;
    input  SCE  ;
    input  SET_B;
    input  VPWR ;
    input  VGND ;
    input  VPB  ;
    input  VNB  ;
    sky130_fd_sc_hvl__sdfstp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .SET_B(SET_B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFSTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxbp: Scan delay flop, non-inverted clock, complementary outputs.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfxbp: Scan delay flop, non-inverted clock, complementary outputs.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__sdfxbp (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q      ;
    wire mux_out    ;
    wire buf0_out_Q ;
    wire not0_out_qn;

    //                                  Delay       Name         Output       Other arguments
    sky130_fd_sc_hvl__udp_mux_2to1                  mux_2to10   (mux_out    , D, SCD, SCE               );
    sky130_fd_sc_hvl__udp_dff$P_pp$PG$N #1 dff0        (buf_Q      , mux_out, CLK, , VPWR, VGND);
    buf                                             buf0        (buf0_out_Q , buf_Q                     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG             pwrgood_pp0 (Q          , buf0_out_Q, VPWR, VGND    );
    not                                             not0        (not0_out_qn, buf_Q                     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG             pwrgood_pp1 (Q_N        , not0_out_qn, VPWR, VGND   );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFXBP_FUNCTIONAL_PP_V


























































































 // FUNCTIONAL




























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFXBP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxbp: Scan delay flop, non-inverted clock, complementary outputs.
 *
 * Verilog wrapper for sdfxbp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__sdfxbp_1 (
    Q   ,
    Q_N ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    output Q_N ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__sdfxbp base (
        .Q(Q),
        .Q_N(Q_N),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/







































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFXBP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxtp: Scan delay flop, non-inverted clock, single output.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdfxtp: Scan delay flop, non-inverted clock, single output.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__sdfxtp (
    Q   ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire buf_Q     ;
    wire mux_out   ;
    wire buf0_out_Q;

    //                                  Delay       Name         Output      Other arguments
    sky130_fd_sc_hvl__udp_mux_2to1                  mux_2to10   (mux_out   , D, SCD, SCE               );
    sky130_fd_sc_hvl__udp_dff$P_pp$PG$N #1 dff0        (buf_Q     , mux_out, CLK, , VPWR, VGND);
    buf                                             buf0        (buf0_out_Q, buf_Q                     );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG             pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND    );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFXTP_FUNCTIONAL_PP_V





















































































 // FUNCTIONAL






















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdfxtp: Scan delay flop, non-inverted clock, single output.
 *
 * Verilog wrapper for sdfxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__sdfxtp_1 (
    Q   ,
    CLK ,
    D   ,
    SCD ,
    SCE ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  CLK ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__sdfxtp base (
        .Q(Q),
        .CLK(CLK),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDFXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdlclkp: Scan gated clock.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdlclkp: Scan gated clock.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__sdlclkp (
    GCLK,
    SCE ,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output GCLK;
    input  SCE ;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire m0      ;
    wire m0n     ;
    wire clkn    ;
    wire SCE_GATE;
    wire GCLK_b  ;

    //                                     Name         Output    Other arguments
    not                                    not0        (m0n     , m0                          );
    not                                    not1        (clkn    , CLK                         );
    nor                                    nor0        (SCE_GATE, GATE, SCE                   );
    sky130_fd_sc_hvl__udp_dlatch$P_pp$PG$N dlatch0     (m0      , SCE_GATE, clkn, , VPWR, VGND);
    and                                    and0        (GCLK_b  , m0n, CLK                    );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG    pwrgood_pp0 (GCLK    , GCLK_b, VPWR, VGND          );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SDLCLKP_FUNCTIONAL_PP_V






















































































 // FUNCTIONAL



























































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDLCLKP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdlclkp: Scan gated clock.
 *
 * Verilog wrapper for sdlclkp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__sdlclkp_1 (
    GCLK,
    SCE ,
    GATE,
    CLK ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output GCLK;
    input  SCE ;
    input  GATE;
    input  CLK ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__sdlclkp base (
        .GCLK(GCLK),
        .SCE(SCE),
        .GATE(GATE),
        .CLK(CLK),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/

































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDLCLKP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdlxtp: ????.
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * sdlxtp: ????.
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__sdlxtp (
    Q   ,
    D   ,
    SCD ,
    SCE ,
    GATE,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Q   ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  GATE;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire mux_out   ;
    wire buf_Q     ;
    wire buf0_out_Q;

    //                                     Delay       Name         Output      Other arguments
    sky130_fd_sc_hvl__udp_mux_2to1                     mux_2to10   (mux_out   , D, SCD, SCE                );
    sky130_fd_sc_hvl__udp_dlatch$P_pp$PG$N #1 dlatch0     (buf_Q     , mux_out, GATE, , VPWR, VGND);
    buf                                                buf0        (buf0_out_Q, buf_Q                      );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG                pwrgood_pp0 (Q         , buf0_out_Q, VPWR, VGND     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__SDLXTP_FUNCTIONAL_PP_V




















































































 // FUNCTIONAL





















































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDLXTP_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * sdlxtp: ????.
 *
 * Verilog wrapper for sdlxtp with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__sdlxtp_1 (
    Q   ,
    D   ,
    SCD ,
    SCE ,
    GATE,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Q   ;
    input  D   ;
    input  SCD ;
    input  SCE ;
    input  GATE;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__sdlxtp base (
        .Q(Q),
        .D(D),
        .SCD(SCD),
        .SCE(SCE),
        .GATE(GATE),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/




































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__SDLXTP_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor2: 2-input exclusive NOR.
 *
 *        Y = !(A ^ B)
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * xnor2: 2-input exclusive NOR.
 *
 *        Y = !(A ^ B)
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__xnor2 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire xnor0_out_Y      ;
    wire pwrgood_pp0_out_Y;

    //                                  Name         Output             Other arguments
    xnor                                xnor0       (xnor0_out_Y      , A, B                   );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_Y, xnor0_out_Y, VPWR, VGND);
    buf                                 buf0        (Y                , pwrgood_pp0_out_Y      );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__XNOR2_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__XNOR2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xnor2: 2-input exclusive NOR.
 *
 *        Y = !(A ^ B)
 *
 * Verilog wrapper for xnor2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__xnor2_1 (
    Y   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__xnor2 base (
        .Y(Y),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__XNOR2_1_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor2: 2-input exclusive OR.
 *
 *       X = A ^ B
 *
 * Verilog top module.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none




/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/





/**
 * xor2: 2-input exclusive OR.
 *
 *       X = A ^ B
 *
 * Verilog simulation functional model.
 */

`timescale 1ns / 1ps
`default_nettype none

// Import user defined primitives.

`celldefine
module sky130_fd_sc_hvl__xor2 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    // Module ports
    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;

    // Local signals
    wire xor0_out_X       ;
    wire pwrgood_pp0_out_X;

    //                                  Name         Output             Other arguments
    xor                                 xor0        (xor0_out_X       , B, A                  );
    sky130_fd_sc_hvl__udp_pwrgood_pp$PG pwrgood_pp0 (pwrgood_pp0_out_X, xor0_out_X, VPWR, VGND);
    buf                                 buf0        (X                , pwrgood_pp0_out_X     );

endmodule
`endcelldefine

`default_nettype wire
  // SKY130_FD_SC_HVL__XOR2_FUNCTIONAL_PP_V






































































 // FUNCTIONAL































































































































 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__XOR2_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */




/**
 * xor2: 2-input exclusive OR.
 *
 *       X = A ^ B
 *
 * Verilog wrapper for xor2 with size of 1 units.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none



/*********************************************************/

`celldefine
module sky130_fd_sc_hvl__xor2_1 (
    X   ,
    A   ,
    B   ,
    VPWR,
    VGND,
    VPB ,
    VNB
);

    output X   ;
    input  A   ;
    input  B   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
    sky130_fd_sc_hvl__xor2 base (
        .X(X),
        .A(A),
        .B(B),
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPB),
        .VNB(VNB)
    );

endmodule
`endcelldefine

/*********************************************************/






























 // USE_POWER_PINS

`default_nettype wire
  // SKY130_FD_SC_HVL__XOR2_1_V


//--------EOF---------

// OpenRAM SRAM model
// Words: 512
// Word size: 32
// Write size: 8

module sky130_sram_2kbyte_1rw1r_32x512_8(

    vccd1,
    vssd1,

// Port 0: RW
    clk0,csb0,web0,wmask0,addr0,din0,dout0,
// Port 1: R
    clk1,csb1,addr1,dout1
  );

  parameter NUM_WMASKS = 4 ;
  parameter DATA_WIDTH = 32 ;
  parameter ADDR_WIDTH = 9 ;
  parameter RAM_DEPTH = 1 << ADDR_WIDTH;
  // FIXME: This delay is arbitrary.
  parameter DELAY = 3 ;
  parameter VERBOSE = 0 ; //Set to 0 to only display warnings
  parameter T_HOLD = 1 ; //Delay to hold dout value after posedge. Value is arbitrary


    inout vccd1;
    inout vssd1;

  input  clk0; // clock
  input   csb0; // active low chip select
  input  web0; // active low write control
  input [NUM_WMASKS-1:0]   wmask0; // write mask
  input [ADDR_WIDTH-1:0]  addr0;
  input [DATA_WIDTH-1:0]  din0;
  output [DATA_WIDTH-1:0] dout0;
  input  clk1; // clock
  input   csb1; // active low chip select
  input [ADDR_WIDTH-1:0]  addr1;
  output [DATA_WIDTH-1:0] dout1;

  reg  csb0_reg;
  reg  web0_reg;
  reg [NUM_WMASKS-1:0]   wmask0_reg;
  reg [ADDR_WIDTH-1:0]  addr0_reg;
  reg [DATA_WIDTH-1:0]  din0_reg;
  reg [DATA_WIDTH-1:0]  dout0;

  reg [DATA_WIDTH-1:0]    mem [0:RAM_DEPTH-1];

  // All inputs are registers
  always @(posedge clk0)
  begin
    csb0_reg = csb0;
    web0_reg = web0;
    wmask0_reg = wmask0;
    addr0_reg = addr0;
    din0_reg = din0;
    #(T_HOLD) dout0 = 32'bx;
    if ( !csb0_reg && web0_reg && VERBOSE ) 
      $display($time," Reading %m addr0=%b dout0=%b",addr0_reg,mem[addr0_reg]);
    if ( !csb0_reg && !web0_reg && VERBOSE )
      $display($time," Writing %m addr0=%b din0=%b wmask0=%b",addr0_reg,din0_reg,wmask0_reg);
  end

  reg  csb1_reg;
  reg [ADDR_WIDTH-1:0]  addr1_reg;
  reg [DATA_WIDTH-1:0]  dout1;

  // All inputs are registers
  always @(posedge clk1)
  begin
    csb1_reg = csb1;
    addr1_reg = addr1;
    if (!csb0 && !web0 && !csb1 && (addr0 == addr1))
         $display($time," WARNING: Writing and reading addr0=%b and addr1=%b simultaneously!",addr0,addr1);
    #(T_HOLD) dout1 = 32'bx;
    if ( !csb1_reg && VERBOSE ) 
      $display($time," Reading %m addr1=%b dout1=%b",addr1_reg,mem[addr1_reg]);
  end


  // Memory Write Block Port 0
  // Write Operation : When web0 = 0, csb0 = 0
  always @ (negedge clk0)
  begin : MEM_WRITE0
    if ( !csb0_reg && !web0_reg ) begin
        if (wmask0_reg[0])
                mem[addr0_reg][7:0] = din0_reg[7:0];
        if (wmask0_reg[1])
                mem[addr0_reg][15:8] = din0_reg[15:8];
        if (wmask0_reg[2])
                mem[addr0_reg][23:16] = din0_reg[23:16];
        if (wmask0_reg[3])
                mem[addr0_reg][31:24] = din0_reg[31:24];
    end
  end

  // Memory Read Block Port 0
  // Read Operation : When web0 = 1, csb0 = 0
  always @ (negedge clk0)
  begin : MEM_READ0
    if (!csb0_reg && web0_reg)
       dout0 <= #(DELAY) mem[addr0_reg];
  end

  // Memory Read Block Port 1
  // Read Operation : When web1 = 1, csb1 = 0
  always @ (negedge clk1)
  begin : MEM_READ1
    if (!csb1_reg)
       dout1 <= #(DELAY) mem[addr1_reg];
  end

endmodule
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

















































 // __GLOBAL_DEFINE_H
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
		parameter BITS = 32
	) (
	
		inout vdda1,	// User area 1 3.3V supply
		inout vdda2,	// User area 2 3.3V supply
		inout vssa1,	// User area 1 analog ground
		inout vssa2,	// User area 2 analog ground
		inout vccd1,	// User area 1 1.8V supply
		inout vccd2,	// User area 2 1.8v supply
		inout vssd1,	// User area 1 digital ground
		inout vssd2,	// User area 2 digital ground
	

		// Wishbone Slave ports (WB MI A)
		input wb_clk_i,
		input wb_rst_i,
		input wbs_stb_i,
		input wbs_cyc_i,
		input wbs_we_i,
		input [3:0] wbs_sel_i,
		input [31:0] wbs_dat_i,
		input [31:0] wbs_adr_i,
		output wbs_ack_o,
		output [31:0] wbs_dat_o,

		// Logic Analyzer Signals
		input  [127:0] la_data_in,
		output [127:0] la_data_out,
		input  [127:0] la_oenb,

		// IOs
		input  [(19 + 19)-1:0] io_in,
		output [(19 + 19)-1:0] io_out,
		output [(19 + 19)-1:0] io_oeb,

		// Analog (direct connection to GPIO pad---use with caution)
		// Note that analog I/O is not available on the 7 lowest-numbered
		// GPIO pads, and so the analog_io indexing is offset from the
		// GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
		inout [(19 + 19)-10:0] analog_io,

		// Independent clock (on independent integer divider)
		input   user_clock2,

		// User maskable interrupt signals
		output [2:0] user_irq
	);

	/*--------------------------------------*/
	/* User project is instantiated  here   */
	/*--------------------------------------*/

	// Caravel wishbone master
	wire caravel_wb_cyc_o;
	wire caravel_wb_stb_o;
	wire caravel_wb_we_o;
	wire[3:0] caravel_wb_sel_o;
	wire[31:0] caravel_wb_data_o;
	wire[27:0] caravel_wb_adr_o;
	wire caravel_wb_ack_i;
	wire caravel_wb_stall_i;
	wire caravel_wb_error_i;
	wire[31:0] caravel_wb_data_i;

	// Caravel
	wire caravel_uart_rx;
	wire caravel_uart_tx;
	wire[3:0] caravel_irq;

	assign user_irq = caravel_irq[2:0];

	// Configuration
	wire[7:0] core0Index;
	wire[7:0] core1Index;
	wire[10:0] manufacturerID;
	wire[15:0] partID;
	wire[3:0] versionID;

	// Debug
	//wire[97:0] soc_probe_in;
	wire[97:0] soc_probe_out;

	ExperiarSoC experiarSoC(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

    	.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.caravel_wb_cyc_o(caravel_wb_cyc_o),
		.caravel_wb_stb_o(caravel_wb_stb_o),
		.caravel_wb_we_o(caravel_wb_we_o),
		.caravel_wb_sel_o(caravel_wb_sel_o),
		.caravel_wb_data_o(caravel_wb_data_o),
		.caravel_wb_adr_o(caravel_wb_adr_o),
		.caravel_wb_ack_i(caravel_wb_ack_i),
		.caravel_wb_stall_i(caravel_wb_stall_i),
		.caravel_wb_error_i(caravel_wb_error_i),
		.caravel_wb_data_i(caravel_wb_data_i),
		.io_in(io_in),
		.io_out(io_out),
		.io_oeb(io_oeb),
		.caravel_uart_rx(caravel_uart_rx),
		.caravel_uart_tx(caravel_uart_tx),
		.caravel_irq(caravel_irq),
		//.probe_in(soc_probe_in),
		.probe_out(soc_probe_out),
		.core0Index(core0Index),
		.core1Index(core1Index),
		.manufacturerID(manufacturerID),
		.partID(partID),
		.versionID(versionID));

	CaravelHost caravelHost(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.wb_clk_i(wb_clk_i),
    	.wb_rst_i(wb_rst_i),
		.wbs_stb_i(wbs_stb_i),
		.wbs_cyc_i(wbs_cyc_i),
		.wbs_we_i(wbs_we_i),
		.wbs_sel_i(wbs_sel_i),
		.wbs_data_i(wbs_dat_i),
		.wbs_adr_i(wbs_adr_i),
		.wbs_ack_o(wbs_ack_o),
		.wbs_data_o(wbs_dat_o),
		.caravel_wb_cyc_o(caravel_wb_cyc_o),
		.caravel_wb_stb_o(caravel_wb_stb_o),
		.caravel_wb_we_o(caravel_wb_we_o),
		.caravel_wb_sel_o(caravel_wb_sel_o),
		.caravel_wb_data_o(caravel_wb_data_o),
		.caravel_wb_adr_o(caravel_wb_adr_o),
		.caravel_wb_ack_i(caravel_wb_ack_i),
		.caravel_wb_stall_i(caravel_wb_stall_i),
		.caravel_wb_error_i(caravel_wb_error_i),
		.caravel_wb_data_i(caravel_wb_data_i),
		// Swap Tx and Rx pins, as these are with reference to the interface
		.caravel_uart_rx(caravel_uart_tx),
		.caravel_uart_tx(caravel_uart_rx),
		.caravel_irq(caravel_irq),
		//.la_data_in(la_data_in),
		.la_data_out(la_data_out),
		//.la_oenb(la_oenb),
		//.probe_in(soc_probe_in),
		.probe_out(soc_probe_out),
		.core0Index(core0Index),
		.core1Index(core1Index),
		.manufacturerID(manufacturerID),
		.partID(partID),
		.versionID(versionID));

	// Add dumby module for art
	Art art(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1)	// User area 1 digital ground

		);

endmodule	// user_project_wrapper

`default_nettype wire
module ExperiarSoC (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		input wire wb_clk_i,
		input wire wb_rst_i,

		// Caravel wishbone master
		input wire caravel_wb_cyc_o,
		input wire caravel_wb_stb_o,
		input wire caravel_wb_we_o,
		input wire[3:0] caravel_wb_sel_o,
		input wire[31:0] caravel_wb_data_o,
		input wire[27:0] caravel_wb_adr_o,
		output wire caravel_wb_ack_i,
		output wire caravel_wb_stall_i,
		output wire caravel_wb_error_i,
		output wire[31:0] caravel_wb_data_i,

		// IOs
		input  wire[(19 + 19)-1:0] io_in,
		output wire[(19 + 19)-1:0] io_out,
		output wire[(19 + 19)-1:0] io_oeb,
		
		// Caravel
		input wire caravel_uart_rx,
		output wire caravel_uart_tx,
		input wire[3:0] caravel_irq,

		// Logic Analyzer Signals
		//input wire[127:0] probe_in,
		output wire[97:0] probe_out,

		// Configuration constants
		input wire[7:0] core0Index,
		input wire[7:0] core1Index,
		input wire[10:0] manufacturerID,
		input wire[15:0] partID,
		input wire[3:0] versionID
	);
	
	localparam SRAM_ADDRESS_SIZE = 9;
	
	// JTAG
	wire jtag_tck;
	wire jtag_tms;
	wire jtag_tdi;
	wire jtag_tdo;

	// Flash
	wire flash_csb;
	wire flash_sck;
	wire flash_io0_we;
	wire flash_io0_write;
	wire flash_io0_read;
	wire flash_io1_we;
	wire flash_io1_write;
	wire flash_io1_read;

	// IRQ
	// wire irq_en;
	// wire irq_in;
	wire[15:0] irq;

	// Wishbone wires
	// Master 0: Caravel

	// Master 1: Core 0
	wire core0_wb_cyc_o;
	wire core0_wb_stb_o;
	wire core0_wb_we_o;
	wire[3:0] core0_wb_sel_o;
	wire[31:0] core0_wb_data_o;
	wire[27:0] core0_wb_adr_o;
	wire core0_wb_ack_i;
	wire core0_wb_stall_i;
	wire core0_wb_error_i;
	wire[31:0] core0_wb_data_i;

	// Master 2: Core 1
	wire core1_wb_cyc_o;
	wire core1_wb_stb_o;
	wire core1_wb_we_o;
	wire[3:0] core1_wb_sel_o;
	wire[31:0] core1_wb_data_o;
	wire[27:0] core1_wb_adr_o;
	wire core1_wb_ack_i;
	wire core1_wb_stall_i;
	wire core1_wb_error_i;
	wire[31:0] core1_wb_data_i;

	// Master 3: dma
	// wire dma_wb_cyc_o = 1'b0;
	// wire dma_wb_stb_o = 1'b0;
	// wire dma_wb_we_o = 1'b0;
	// wire[3:0] dma_wb_sel_o = 4'b0;
	// wire[31:0] dma_wb_data_o = 32'b0;
	// wire[27:0] dma_wb_adr_o = 28'b0;
	// wire dma_wb_ack_i;
	// wire dma_wb_stall_i;
	// wire dma_wb_error_i;
	// wire[31:0] dma_wb_data_i;

	// Slave 0
	wire core0Memory_wb_cyc_i;
	wire core0Memory_wb_stb_i;
	wire core0Memory_wb_we_i;
	wire[3:0] core0Memory_wb_sel_i;
	wire[31:0] core0Memory_wb_data_i;
	wire[23:0] core0Memory_wb_adr_i;
	wire core0Memory_wb_ack_o;
	wire core0Memory_wb_stall_o;
	wire core0Memory_wb_error_o;
	wire[31:0] core0Memory_wb_data_o;

	// Slave 1
	wire core1Memory_wb_cyc_i;
	wire core1Memory_wb_stb_i;
	wire core1Memory_wb_we_i;
	wire[3:0] core1Memory_wb_sel_i;
	wire[31:0] core1Memory_wb_data_i;
	wire[23:0] core1Memory_wb_adr_i;
	wire core1Memory_wb_ack_o;
	wire core1Memory_wb_stall_o;
	wire core1Memory_wb_error_o;
	wire[31:0] core1Memory_wb_data_o;

	// Slave 2
	wire videoMemory_wb_cyc_i;
	wire videoMemory_wb_stb_i;
	wire videoMemory_wb_we_i;
	wire[3:0] videoMemory_wb_sel_i;
	wire[31:0] videoMemory_wb_data_i;
	wire[23:0] videoMemory_wb_adr_i;
	wire videoMemory_wb_ack_o;
	wire videoMemory_wb_stall_o;
	wire videoMemory_wb_error_o;
	wire[31:0] videoMemory_wb_data_o;

	// Slave 3
	wire peripherals_wb_cyc_i;
	wire peripherals_wb_stb_i;
	wire peripherals_wb_we_i;
	wire[3:0] peripherals_wb_sel_i;
	wire[31:0] peripherals_wb_data_i;
	wire[23:0] peripherals_wb_adr_i;
	wire peripherals_wb_ack_o;
	wire peripherals_wb_stall_o;
	wire peripherals_wb_error_o;
	wire[31:0] peripherals_wb_data_o;

	// Slave 4
	wire flash_wb_cyc_i;
	wire flash_wb_stb_i;
	wire flash_wb_we_i;
	wire[3:0] flash_wb_sel_i;
	wire[31:0] flash_wb_data_i;
	wire[23:0] flash_wb_adr_i;
	wire flash_wb_ack_o;
	wire flash_wb_stall_o;
	wire flash_wb_error_o;
	wire[31:0] flash_wb_data_o;

	// wire[2:0] probe_master0_currentSlave;
	// wire[2:0] probe_master1_currentSlave;
	// wire[2:0] probe_master2_currentSlave;
	// wire[2:0] probe_master3_currentSlave;
	// wire[1:0] probe_slave0_currentMaster;
	// wire[1:0] probe_slave1_currentMaster;
	// wire[1:0] probe_slave2_currentMaster;
	// wire[1:0] probe_slave3_currentMaster;
	// wire[1:0] probe_slave4_currentMaster;

	// wire[15:0] probe_wishboneInterconnect = {
	// 	probe_slave3_currentMaster,
	// 	probe_slave2_currentMaster,
	// 	probe_slave1_currentMaster,
	// 	probe_slave0_currentMaster,
	// 	probe_master3_currentSlave[1:0],
	// 	probe_master2_currentSlave[1:0],
	// 	probe_master1_currentSlave[1:0],
	// 	probe_master0_currentSlave[1:0]
	// };

	wire[1:0] probe_master0_currentSlave;
	wire[1:0] probe_master1_currentSlave;
	wire[1:0] probe_master2_currentSlave;
	wire[1:0] probe_master3_currentSlave;
	wire[1:0] probe_slave0_currentMaster;
	wire[1:0] probe_slave1_currentMaster;
	wire[1:0] probe_slave2_currentMaster;
	wire[1:0] probe_slave3_currentMaster;

	wire[15:0] probe_wishboneInterconnect = {
		probe_slave3_currentMaster,
		probe_slave2_currentMaster,
		probe_slave1_currentMaster,
		probe_slave0_currentMaster,
		probe_master3_currentSlave,
		probe_master2_currentSlave,
		probe_master1_currentSlave,
		probe_master0_currentSlave
	};

	//-------------------------------------------------//
	//---------------------Wishbone--------------------//
	//-------------------------------------------------//

	WishboneInterconnect wishboneInterconnect(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.master0_wb_cyc_o(caravel_wb_cyc_o),
		.master0_wb_stb_o(caravel_wb_stb_o),
		.master0_wb_we_o(caravel_wb_we_o),
		.master0_wb_sel_o(caravel_wb_sel_o),
		.master0_wb_data_o(caravel_wb_data_o),
		.master0_wb_adr_o(caravel_wb_adr_o),
		.master0_wb_ack_i(caravel_wb_ack_i),
		.master0_wb_stall_i(caravel_wb_stall_i),
		.master0_wb_error_i(caravel_wb_error_i),
		.master0_wb_data_i(caravel_wb_data_i),
		.master1_wb_cyc_o(core0_wb_cyc_o),
		.master1_wb_stb_o(core0_wb_stb_o),
		.master1_wb_we_o(core0_wb_we_o),
		.master1_wb_sel_o(core0_wb_sel_o),
		.master1_wb_data_o(core0_wb_data_o),
		.master1_wb_adr_o(core0_wb_adr_o),
		.master1_wb_ack_i(core0_wb_ack_i),
		.master1_wb_stall_i(core0_wb_stall_i),
		.master1_wb_error_i(core0_wb_error_i),
		.master1_wb_data_i(core0_wb_data_i),
		.master2_wb_cyc_o(core1_wb_cyc_o),
		.master2_wb_stb_o(core1_wb_stb_o),
		.master2_wb_we_o(core1_wb_we_o),
		.master2_wb_sel_o(core1_wb_sel_o),
		.master2_wb_data_o(core1_wb_data_o),
		.master2_wb_adr_o(core1_wb_adr_o),
		.master2_wb_ack_i(core1_wb_ack_i),
		.master2_wb_stall_i(core1_wb_stall_i),
		.master2_wb_error_i(core1_wb_error_i),
		.master2_wb_data_i(core1_wb_data_i),
		// .master3_wb_cyc_o(dma_wb_cyc_o),
		// .master3_wb_stb_o(dma_wb_stb_o),
		// .master3_wb_we_o(dma_wb_we_o),
		// .master3_wb_sel_o(dma_wb_sel_o),
		// .master3_wb_data_o(dma_wb_data_o),
		// .master3_wb_adr_o(dma_wb_adr_o),
		// .master3_wb_ack_i(dma_wb_ack_i),
		// .master3_wb_stall_i(dma_wb_stall_i),
		// .master3_wb_error_i(dma_wb_error_i),
		// .master3_wb_data_i(dma_wb_data_i),
		.slave0_wb_cyc_i(core0Memory_wb_cyc_i),
		.slave0_wb_stb_i(core0Memory_wb_stb_i),
		.slave0_wb_we_i(core0Memory_wb_we_i),
		.slave0_wb_sel_i(core0Memory_wb_sel_i),
		.slave0_wb_data_i(core0Memory_wb_data_i),
		.slave0_wb_adr_i(core0Memory_wb_adr_i),
		.slave0_wb_ack_o(core0Memory_wb_ack_o),
		.slave0_wb_stall_o(core0Memory_wb_stall_o),
		.slave0_wb_error_o(core0Memory_wb_error_o),
		.slave0_wb_data_o(core0Memory_wb_data_o),
		.slave1_wb_cyc_i(core1Memory_wb_cyc_i),
		.slave1_wb_stb_i(core1Memory_wb_stb_i),
		.slave1_wb_we_i(core1Memory_wb_we_i),
		.slave1_wb_sel_i(core1Memory_wb_sel_i),
		.slave1_wb_data_i(core1Memory_wb_data_i),
		.slave1_wb_adr_i(core1Memory_wb_adr_i),
		.slave1_wb_ack_o(core1Memory_wb_ack_o),
		.slave1_wb_stall_o(core1Memory_wb_stall_o),
		.slave1_wb_error_o(core1Memory_wb_error_o),
		.slave1_wb_data_o(core1Memory_wb_data_o),
		.slave2_wb_cyc_i(videoMemory_wb_cyc_i),
		.slave2_wb_stb_i(videoMemory_wb_stb_i),
		.slave2_wb_we_i(videoMemory_wb_we_i),
		.slave2_wb_sel_i(videoMemory_wb_sel_i),
		.slave2_wb_data_i(videoMemory_wb_data_i),
		.slave2_wb_adr_i(videoMemory_wb_adr_i),
		.slave2_wb_ack_o(videoMemory_wb_ack_o),
		.slave2_wb_stall_o(videoMemory_wb_stall_o),
		.slave2_wb_error_o(videoMemory_wb_error_o),
		.slave2_wb_data_o(videoMemory_wb_data_o),
		.slave3_wb_cyc_i(peripherals_wb_cyc_i),
		.slave3_wb_stb_i(peripherals_wb_stb_i),
		.slave3_wb_we_i(peripherals_wb_we_i),
		.slave3_wb_sel_i(peripherals_wb_sel_i),
		.slave3_wb_data_i(peripherals_wb_data_i),
		.slave3_wb_adr_i(peripherals_wb_adr_i),
		.slave3_wb_ack_o(peripherals_wb_ack_o),
		.slave3_wb_stall_o(peripherals_wb_stall_o),
		.slave3_wb_error_o(peripherals_wb_error_o),
		.slave3_wb_data_o(peripherals_wb_data_o),
		.slave4_wb_cyc_i(flash_wb_cyc_i),
		.slave4_wb_stb_i(flash_wb_stb_i),
		.slave4_wb_we_i(flash_wb_we_i),
		.slave4_wb_sel_i(flash_wb_sel_i),
		.slave4_wb_data_i(flash_wb_data_i),
		.slave4_wb_adr_i(flash_wb_adr_i),
		.slave4_wb_ack_o(flash_wb_ack_o),
		.slave4_wb_stall_o(flash_wb_stall_o),
		.slave4_wb_error_o(flash_wb_error_o),
		.slave4_wb_data_o(flash_wb_data_o),
		.probe_master0_currentSlave(probe_master0_currentSlave),
		.probe_master1_currentSlave(probe_master1_currentSlave),
		.probe_master2_currentSlave(probe_master2_currentSlave),
		.probe_master3_currentSlave(probe_master3_currentSlave),
		.probe_slave0_currentMaster(probe_slave0_currentMaster),
		.probe_slave1_currentMaster(probe_slave1_currentMaster),
		.probe_slave2_currentMaster(probe_slave2_currentMaster),
		.probe_slave3_currentMaster(probe_slave3_currentMaster));//,
		//.probe_slave4_currentMaster(probe_slave4_currentMaster));

	//-------------------------------------------------//
	//----------------------CORE0----------------------//
	//-------------------------------------------------//
	
	// JTAG interface
	wire core0_tdi;
	wire core0_tdo;

	// SRAM rw port
	wire core0SRAM_clk0;
	wire[1:0] core0SRAM_csb0;
	wire core0SRAM_web0;
	wire[3:0] core0SRAM_wmask0;
	wire[SRAM_ADDRESS_SIZE-1:0] core0SRAM_addr0;
	wire[31:0] core0SRAM_din0;
	wire[63:0] core0SRAM_dout0;

	// SRAM r port
	wire core0SRAM_clk1;
	wire[1:0] core0SRAM_csb1;
	wire[SRAM_ADDRESS_SIZE-1:0] core0SRAM_addr1;
	wire[63:0] core0SRAM_dout1;

	// Logic probes
	wire probe_core0_state;
	wire[1:0] probe_core0_env;
	wire[31:0] probe_core0_programCounter;
	wire[4:0] probe_core0_jtagInstruction;

	wire[39:0] probe_core0 = {
		probe_core0_state,
		probe_core0_env,
		probe_core0_programCounter,
		probe_core0_jtagInstruction
	};

	ExperiarCore core0 (

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.coreIndex(core0Index),
		.manufacturerID(manufacturerID),
		.partID(partID),
		.versionID(versionID),
		.jtag_tck(jtag_tck),
		.jtag_tms(jtag_tms),
		.jtag_tdi(core0_tdi),
		.jtag_tdo(core0_tdo),
		.irq(irq),
		.core_wb_cyc_o(core0_wb_cyc_o),
		.core_wb_stb_o(core0_wb_stb_o),
		.core_wb_we_o(core0_wb_we_o),
		.core_wb_sel_o(core0_wb_sel_o),
		.core_wb_data_o(core0_wb_data_o),
		.core_wb_adr_o(core0_wb_adr_o),
		.core_wb_ack_i(core0_wb_ack_i),
		.core_wb_stall_i(core0_wb_stall_i),
		.core_wb_error_i(core0_wb_error_i),
		.core_wb_data_i(core0_wb_data_i),
		.localMemory_wb_cyc_i(core0Memory_wb_cyc_i),
		.localMemory_wb_stb_i(core0Memory_wb_stb_i),
		.localMemory_wb_we_i(core0Memory_wb_we_i),
		.localMemory_wb_sel_i(core0Memory_wb_sel_i),
		.localMemory_wb_data_i(core0Memory_wb_data_i),
		.localMemory_wb_adr_i(core0Memory_wb_adr_i),
		.localMemory_wb_ack_o(core0Memory_wb_ack_o),
		.localMemory_wb_stall_o(core0Memory_wb_stall_o),
		.localMemory_wb_error_o(core0Memory_wb_error_o),
		.localMemory_wb_data_o(core0Memory_wb_data_o),
		.clk0(core0SRAM_clk0),
		.csb0(core0SRAM_csb0),
		.web0(core0SRAM_web0),
		.wmask0(core0SRAM_wmask0),
		.addr0(core0SRAM_addr0),
		.din0(core0SRAM_din0),
		.dout0(core0SRAM_dout0),
		.clk1(core0SRAM_clk1),
		.csb1(core0SRAM_csb1),
		.addr1(core0SRAM_addr1),
		.dout1(core0SRAM_dout1),
		.probe_state(probe_core0_state),
		.probe_env(probe_core0_env),
		.probe_programCounter(probe_core0_programCounter),
		.probe_jtagInstruction(probe_core0_jtagInstruction));

	wire[31:0] core0SRAM0_dout0;
	wire[31:0] core0SRAM0_dout1;
	sky130_sram_2kbyte_1rw1r_32x512_8 core0SRAM0(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(core0SRAM_clk0),
		.csb0(core0SRAM_csb0[0]),
		.web0(core0SRAM_web0),
		.wmask0(core0SRAM_wmask0),
		.addr0(core0SRAM_addr0),
		.din0(core0SRAM_din0),
		.dout0(core0SRAM0_dout0),
		.clk1(core0SRAM_clk1),
		.csb1(core0SRAM_csb1[0]),
		.addr1(core0SRAM_addr1),
		.dout1(core0SRAM0_dout1));

	wire[31:0] core0SRAM1_dout0;
	wire[31:0] core0SRAM1_dout1;
	sky130_sram_2kbyte_1rw1r_32x512_8 core0SRAM1(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(core0SRAM_clk0),
		.csb0(core0SRAM_csb0[1]),
		.web0(core0SRAM_web0),
		.wmask0(core0SRAM_wmask0),
		.addr0(core0SRAM_addr0),
		.din0(core0SRAM_din0),
		.dout0(core0SRAM1_dout0),
		.clk1(core0SRAM_clk1),
		.csb1(core0SRAM_csb1[1]),
		.addr1(core0SRAM_addr1),
		.dout1(core0SRAM1_dout1));

	assign core0SRAM_dout0 = { core0SRAM1_dout0, core0SRAM0_dout0 };
	assign core0SRAM_dout1 = { core0SRAM1_dout1, core0SRAM0_dout1 };

	//-------------------------------------------------//
	//----------------------CORE1----------------------//
	//-------------------------------------------------//
	
	// JTAG interface
	wire core1_tdi;
	wire core1_tdo;
	
	// SRAM rw port
	wire core1SRAM_clk0;
	wire[1:0] core1SRAM_csb0;
	wire core1SRAM_web0;
	wire[3:0] core1SRAM_wmask0;
	wire[SRAM_ADDRESS_SIZE-1:0] core1SRAM_addr0;
	wire[31:0] core1SRAM_din0;
	wire[63:0] core1SRAM_dout0;

	// SRAM r port
	wire core1SRAM_clk1;
	wire[1:0] core1SRAM_csb1;
	wire[SRAM_ADDRESS_SIZE-1:0] core1SRAM_addr1;
	wire[63:0] core1SRAM_dout1;

	// Logic probes
	wire probe_core1_state;
	wire[1:0] probe_core1_env;
	wire[31:0] probe_core1_programCounter;
	wire[4:0] probe_core1_jtagInstruction;

	wire[39:0] probe_core1 = {
		probe_core1_state,
		probe_core1_env,
		probe_core1_programCounter,
		probe_core1_jtagInstruction
	};

	ExperiarCore core1 (

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.coreIndex(core1Index),
		.manufacturerID(manufacturerID),
		.partID(partID),
		.versionID(versionID),
		.jtag_tck(jtag_tck),
		.jtag_tms(jtag_tms),
		.jtag_tdi(core1_tdi),
		.jtag_tdo(core1_tdo),
		.irq(irq),
		.core_wb_cyc_o(core1_wb_cyc_o),
		.core_wb_stb_o(core1_wb_stb_o),
		.core_wb_we_o(core1_wb_we_o),
		.core_wb_sel_o(core1_wb_sel_o),
		.core_wb_data_o(core1_wb_data_o),
		.core_wb_adr_o(core1_wb_adr_o),
		.core_wb_ack_i(core1_wb_ack_i),
		.core_wb_stall_i(core1_wb_stall_i),
		.core_wb_error_i(core1_wb_error_i),
		.core_wb_data_i(core1_wb_data_i),
		.localMemory_wb_cyc_i(core1Memory_wb_cyc_i),
		.localMemory_wb_stb_i(core1Memory_wb_stb_i),
		.localMemory_wb_we_i(core1Memory_wb_we_i),
		.localMemory_wb_sel_i(core1Memory_wb_sel_i),
		.localMemory_wb_data_i(core1Memory_wb_data_i),
		.localMemory_wb_adr_i(core1Memory_wb_adr_i),
		.localMemory_wb_ack_o(core1Memory_wb_ack_o),
		.localMemory_wb_stall_o(core1Memory_wb_stall_o),
		.localMemory_wb_error_o(core1Memory_wb_error_o),
		.localMemory_wb_data_o(core1Memory_wb_data_o),
		.clk0(core1SRAM_clk0),
		.csb0(core1SRAM_csb0),
		.web0(core1SRAM_web0),
		.wmask0(core1SRAM_wmask0),
		.addr0(core1SRAM_addr0),
		.din0(core1SRAM_din0),
		.dout0(core1SRAM_dout0),
		.clk1(core1SRAM_clk1),
		.csb1(core1SRAM_csb1),
		.addr1(core1SRAM_addr1),
		.dout1(core1SRAM_dout1),
		.probe_state(probe_core1_state),
		.probe_env(probe_core1_env),
		.probe_programCounter(probe_core1_programCounter),
		.probe_jtagInstruction(probe_core1_jtagInstruction));

	wire[31:0] core1SRAM0_dout0;
	wire[31:0] core1SRAM0_dout1;
	sky130_sram_2kbyte_1rw1r_32x512_8 core1SRAM0(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(core1SRAM_clk0),
		.csb0(core1SRAM_csb0[0]),
		.web0(core1SRAM_web0),
		.wmask0(core1SRAM_wmask0),
		.addr0(core1SRAM_addr0),
		.din0(core1SRAM_din0),
		.dout0(core1SRAM0_dout0),
		.clk1(core1SRAM_clk1),
		.csb1(core1SRAM_csb1[0]),
		.addr1(core1SRAM_addr1),
		.dout1(core1SRAM0_dout1));

	wire[31:0] core1SRAM1_dout0;
	wire[31:0] core1SRAM1_dout1;
	sky130_sram_2kbyte_1rw1r_32x512_8 core1SRAM1(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(core1SRAM_clk0),
		.csb0(core1SRAM_csb0[1]),
		.web0(core1SRAM_web0),
		.wmask0(core1SRAM_wmask0),
		.addr0(core1SRAM_addr0),
		.din0(core1SRAM_din0),
		.dout0(core1SRAM1_dout0),
		.clk1(core1SRAM_clk1),
		.csb1(core1SRAM_csb1[1]),
		.addr1(core1SRAM_addr1),
		.dout1(core1SRAM1_dout1));

	assign core1SRAM_dout0 = { core1SRAM1_dout0, core1SRAM0_dout0 };
	assign core1SRAM_dout1 = { core1SRAM1_dout1, core1SRAM0_dout1 };

	//-------------------------------------------------//
	//----------------------Flash----------------------//
	//-------------------------------------------------//

	// Video SRAM rw port
	wire flashSRAM_clk0;
	wire flashSRAM_csb0;
	wire flashSRAM_web0;
	wire[3:0] flashSRAM_wmask0;
	wire[SRAM_ADDRESS_SIZE-1:0] flashSRAM_addr0;
	wire[31:0] flashSRAM_din0;
	wire[31:0] flashSRAM_dout0;

	// Video SRAM r port
	wire flashSRAM_clk1;
	wire flashSRAM_csb1;
	wire[SRAM_ADDRESS_SIZE-1:0] flashSRAM_addr1;
	wire[31:0] flashSRAM_dout1;

	Flash flash(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_stb_i(flash_wb_stb_i),
		.wb_cyc_i(flash_wb_cyc_i),
		.wb_we_i(flash_wb_we_i),
		.wb_sel_i(flash_wb_sel_i),
		.wb_data_i(flash_wb_data_i),
		.wb_adr_i(flash_wb_adr_i),
		.wb_ack_o(flash_wb_ack_o),
		.wb_stall_o(flash_wb_stall_o),
		.wb_error_o(flash_wb_error_o),
		.wb_data_o(flash_wb_data_o),
		.flash_csb(flash_csb),
		.flash_sck(flash_sck),
		.flash_io0_we(flash_io0_we),
		.flash_io0_write(flash_io0_write),
		.flash_io0_read(flash_io0_read),
		.flash_io1_we(flash_io1_we),
		.flash_io1_write(flash_io1_write),
		.flash_io1_read(flash_io1_read),
		.sram_clk0(flashSRAM_clk0),
		.sram_csb0(flashSRAM_csb0),
		.sram_web0(flashSRAM_web0),
		.sram_wmask0(flashSRAM_wmask0),
		.sram_addr0(flashSRAM_addr0),
		.sram_din0(flashSRAM_din0),
		.sram_dout0(flashSRAM_dout0),
		.sram_clk1(flashSRAM_clk1),
		.sram_csb1(flashSRAM_csb1),
		.sram_addr1(flashSRAM_addr1),
		.sram_dout1(flashSRAM_dout1));

		sky130_sram_2kbyte_1rw1r_32x512_8 flashSRAM(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(flashSRAM_clk0),
		.csb0(flashSRAM_csb0),
		.web0(flashSRAM_web0),
		.wmask0(flashSRAM_wmask0),
		.addr0(flashSRAM_addr0),
		.din0(flashSRAM_din0),
		.dout0(flashSRAM_dout0),
		.clk1(flashSRAM_clk1),
		.csb1(flashSRAM_csb1),
		.addr1(flashSRAM_addr1),
		.dout1(flashSRAM_dout1)
	);

	//-------------------------------------------------//
	//----------------------Video----------------------//
	//-------------------------------------------------//

	// VGA
	wire[1:0] vga_r;
	wire[1:0] vga_g;
	wire[1:0] vga_b;
	wire vga_vsync;
	wire vga_hsync;

	// Left Video SRAM rw port
	wire videoSRAMLeft_clk0;
	wire[1:0] videoSRAMLeft_csb0;
	wire videoSRAMLeft_web0;
	wire[3:0] videoSRAMLeft_wmask0;
	wire[SRAM_ADDRESS_SIZE-1:0] videoSRAMLeft_addr0;
	wire[31:0] videoSRAMLeft_din0;
	wire[63:0] videoSRAMLeft_dout0;

	// Left Video SRAM r port
	wire videoSRAMLeft_clk1;
	wire[1:0] videoSRAMLeft_csb1;
	wire[SRAM_ADDRESS_SIZE-1:0] videoSRAMLeft_addr1;
	wire[63:0] videoSRAMLeft_dout1;

	// Right Video SRAM rw port
	wire videoSRAMRight_clk0;
	wire[1:0] videoSRAMRight_csb0;
	wire videoSRAMRight_web0;
	wire[3:0] videoSRAMRight_wmask0;
	wire[SRAM_ADDRESS_SIZE-1:0] videoSRAMRight_addr0;
	wire[31:0] videoSRAMRight_din0;
	wire[63:0] videoSRAMRight_dout0;

	// Right Video SRAM r port
	wire videoSRAMRight_clk1;
	wire[1:0] videoSRAMRight_csb1;
	wire[SRAM_ADDRESS_SIZE-1:0] videoSRAMRight_addr1;
	wire[63:0] videoSRAMRight_dout1;

	wire[1:0] video_irq;
	Video video(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_stb_i(videoMemory_wb_stb_i),
		.wb_cyc_i(videoMemory_wb_cyc_i),
		.wb_we_i(videoMemory_wb_we_i),
		.wb_sel_i(videoMemory_wb_sel_i),
		.wb_data_i(videoMemory_wb_data_i),
		.wb_adr_i(videoMemory_wb_adr_i),
		.wb_ack_o(videoMemory_wb_ack_o),
		.wb_stall_o(videoMemory_wb_stall_o),
		.wb_error_o(videoMemory_wb_error_o),
		.wb_data_o(videoMemory_wb_data_o),
		.video_irq(video_irq),
		.sram0_clk0(videoSRAMLeft_clk0),
		.sram0_csb0(videoSRAMLeft_csb0),
		.sram0_web0(videoSRAMLeft_web0),
		.sram0_wmask0(videoSRAMLeft_wmask0),
		.sram0_addr0(videoSRAMLeft_addr0),
		.sram0_din0(videoSRAMLeft_din0),
		.sram0_dout0(videoSRAMLeft_dout0),
		.sram0_clk1(videoSRAMLeft_clk1),
		.sram0_csb1(videoSRAMLeft_csb1),
		.sram0_addr1(videoSRAMLeft_addr1),
		.sram0_dout1(videoSRAMLeft_dout1),
		.sram1_clk0(videoSRAMRight_clk0),
		.sram1_csb0(videoSRAMRight_csb0),
		.sram1_web0(videoSRAMRight_web0),
		.sram1_wmask0(videoSRAMRight_wmask0),
		.sram1_addr0(videoSRAMRight_addr0),
		.sram1_din0(videoSRAMRight_din0),
		.sram1_dout0(videoSRAMRight_dout0),
		.sram1_clk1(videoSRAMRight_clk1),
		.sram1_csb1(videoSRAMRight_csb1),
		.sram1_addr1(videoSRAMRight_addr1),
		.sram1_dout1(videoSRAMRight_dout1),
		//.vga_clk(wb_clk_i),
		.vga_r(vga_r),
		.vga_g(vga_g),
		.vga_b(vga_b),
		.vga_vsync(vga_vsync),
		.vga_hsync(vga_hsync));

	wire[31:0] videoSRAM0_dout0;
	wire[31:0] videoSRAM0_dout1;
	sky130_sram_2kbyte_1rw1r_32x512_8 videoSRAM0(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(videoSRAMLeft_clk0),
		.csb0(videoSRAMLeft_csb0[0]),
		.web0(videoSRAMLeft_web0),
		.wmask0(videoSRAMLeft_wmask0),
		.addr0(videoSRAMLeft_addr0),
		.din0(videoSRAMLeft_din0),
		.dout0(videoSRAM0_dout0),
		.clk1(videoSRAMLeft_clk1),
		.csb1(videoSRAMLeft_csb1[0]),
		.addr1(videoSRAMLeft_addr1),
		.dout1(videoSRAM0_dout1)
	);

	wire[31:0] videoSRAM1_dout0;
	wire[31:0] videoSRAM1_dout1;
	sky130_sram_2kbyte_1rw1r_32x512_8 videoSRAM1(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(videoSRAMLeft_clk0),
		.csb0(videoSRAMLeft_csb0[1]),
		.web0(videoSRAMLeft_web0),
		.wmask0(videoSRAMLeft_wmask0),
		.addr0(videoSRAMLeft_addr0),
		.din0(videoSRAMLeft_din0),
		.dout0(videoSRAM1_dout0),
		.clk1(videoSRAMLeft_clk1),
		.csb1(videoSRAMLeft_csb1[1]),
		.addr1(videoSRAMLeft_addr1),
		.dout1(videoSRAM1_dout1)
	);

	assign videoSRAMLeft_dout0 = { videoSRAM1_dout0, videoSRAM0_dout0 };
	assign videoSRAMLeft_dout1 = { videoSRAM1_dout1, videoSRAM0_dout1 };

	wire[31:0] videoSRAM2_dout0;
	wire[31:0] videoSRAM2_dout1;
	sky130_sram_2kbyte_1rw1r_32x512_8 videoSRAM2(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(videoSRAMRight_clk0),
		.csb0(videoSRAMRight_csb0[0]),
		.web0(videoSRAMRight_web0),
		.wmask0(videoSRAMRight_wmask0),
		.addr0(videoSRAMRight_addr0),
		.din0(videoSRAMRight_din0),
		.dout0(videoSRAM2_dout0),
		.clk1(videoSRAMRight_clk1),
		.csb1(videoSRAMRight_csb1[0]),
		.addr1(videoSRAMRight_addr1),
		.dout1(videoSRAM2_dout1)
	);

	wire[31:0] videoSRAM3_dout0;
	wire[31:0] videoSRAM3_dout1;
	sky130_sram_2kbyte_1rw1r_32x512_8 videoSRAM3(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk0(videoSRAMRight_clk0),
		.csb0(videoSRAMRight_csb0[1]),
		.web0(videoSRAMRight_web0),
		.wmask0(videoSRAMRight_wmask0),
		.addr0(videoSRAMRight_addr0),
		.din0(videoSRAMRight_din0),
		.dout0(videoSRAM3_dout0),
		.clk1(videoSRAMRight_clk1),
		.csb1(videoSRAMRight_csb1[1]),
		.addr1(videoSRAMRight_addr1),
		.dout1(videoSRAM3_dout1)
	);

	assign videoSRAMRight_dout0 = { videoSRAM3_dout0, videoSRAM2_dout0 };
	assign videoSRAMRight_dout1 = { videoSRAM3_dout1, videoSRAM2_dout1 };

	//-------------------------------------------------//
	//-------------------Peripherals-------------------//
	//-------------------------------------------------//
	wire[1:0] probe_blink;
	wire[9:0] peripheral_irq;
	Peripherals peripherals(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_stb_i(peripherals_wb_stb_i),
		.wb_cyc_i(peripherals_wb_cyc_i),
		.wb_we_i(peripherals_wb_we_i),
		.wb_sel_i(peripherals_wb_sel_i),
		.wb_data_i(peripherals_wb_data_i),
		.wb_adr_i(peripherals_wb_adr_i),
		.wb_ack_o(peripherals_wb_ack_o),
		.wb_stall_o(peripherals_wb_stall_o),
		.wb_error_o(peripherals_wb_error_o),
		.wb_data_o(peripherals_wb_data_o),
		.io_in(io_in),
		.io_out(io_out),
		.io_oeb(io_oeb),
		.internal_uart_rx(caravel_uart_rx),
		.internal_uart_tx(caravel_uart_tx),
		.jtag_tck(jtag_tck),
		.jtag_tms(jtag_tms),
		.jtag_tdi(jtag_tdi),
		.jtag_tdo(jtag_tdo),
		.flash_csb(flash_csb),
		.flash_sck(flash_sck),
		.flash_io0_we(flash_io0_we),
		.flash_io0_write(flash_io0_write),
		.flash_io0_read(flash_io0_read),
		.flash_io1_we(flash_io1_we),
		.flash_io1_write(flash_io1_write),
		.flash_io1_read(flash_io1_read),
		//.irq_en(irq_en),
		//.irq_in(irq_in),
		.peripheral_irq(peripheral_irq),
		.vga_r(vga_r),
		.vga_g(vga_g),
		.vga_b(vga_b),
		.vga_vsync(vga_vsync),
		.vga_hsync(vga_hsync),
		.probe_blink(probe_blink));

	//-------------------------------------------------//
	//-----------------------DMA-----------------------//
	//-------------------------------------------------//

	//DMA dma();

	assign core0_tdi = jtag_tdi;
	assign core1_tdi = core0_tdo;
	assign jtag_tdo = core1_tdo;

	assign probe_out = {
		probe_core1,				// 40
		probe_core0,				// 40
		probe_wishboneInterconnect,	// 16
		probe_blink					// 2
	};

	//-------------------------------------------------//
	//-----------------------IRQ-----------------------//
	//-------------------------------------------------//

	assign irq = { caravel_irq, video_irq, peripheral_irq };

endmodulemodule CaravelHost (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground

		input wire wb_clk_i,
		input wire wb_rst_i,

		// Wishbone Slave port from caravel
		input wbs_stb_i,
		input wbs_cyc_i,
		input wbs_we_i,
		input [3:0] wbs_sel_i,
		input [31:0] wbs_data_i,
		input [31:0] wbs_adr_i,
		output wbs_ack_o,
		output [31:0] wbs_data_o,

		// Caravel wishbone master
		output wire caravel_wb_cyc_o,
		output wire caravel_wb_stb_o,
		output wire caravel_wb_we_o,
		output wire[3:0] caravel_wb_sel_o,
		output wire[31:0] caravel_wb_data_o,
		output wire[27:0] caravel_wb_adr_o,
		input wire caravel_wb_ack_i,
		input wire caravel_wb_stall_i,
		input wire caravel_wb_error_i,
		input wire[31:0] caravel_wb_data_i,
		
		// Caravel UART
		input wire caravel_uart_rx,
		output wire caravel_uart_tx,

		// Caravel IRQ
		output wire[3:0] caravel_irq,

		// Logic probes
		// input wire[127:0] la_data_in,
		output wire[127:0] la_data_out,
		// input wire[127:0] la_oenb,

		//output wire[127:0] probe_in,
		input wire[97:0] probe_out,

		// Configuration constants
		output wire[7:0] core0Index,
		output wire[7:0] core1Index,
		output wire[10:0] manufacturerID,
		output wire[15:0] partID,
		output wire[3:0] versionID
	);

	localparam USER_SPACE_ADDRESS = 4'h3;
	localparam HOST_PERIPHERAL_ADDRESS = 4'hF;

	assign core0Index = 8'h00;
	assign core1Index = 8'h01;
	assign manufacturerID = 11'h000;
	assign partID = 16'hCD55;
	assign versionID = 4'h0;

	wire userSpace_wb_cyc_i;
	wire userSpace_wb_stb_i;
	wire userSpace_wb_we_i;
	wire[3:0] userSpace_wb_sel_i;
	wire[31:0] userSpace_wb_data_i;
	wire[31:0] userSpace_wb_adr_i;
	reg userSpace_wb_ack_o;
	wire[31:0] userSpace_wb_data_o;

	WBAddressExtension wbAddressExtension(
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wbs_cyc_i(wbs_cyc_i),
		.wbs_stb_i(wbs_stb_i),
		.wbs_we_i(wbs_we_i),
		.wbs_sel_i(wbs_sel_i),
		.wbs_adr_i(wbs_adr_i),
		.wbs_data_i(wbs_data_i),
		.wbs_ack_o(wbs_ack_o),
		.wbs_data_o(wbs_data_o),
		.userSpace_wb_cyc_i(userSpace_wb_cyc_i),
		.userSpace_wb_stb_i(userSpace_wb_stb_i),
		.userSpace_wb_we_i(userSpace_wb_we_i),
		.userSpace_wb_sel_i(userSpace_wb_sel_i),
		.userSpace_wb_adr_i(userSpace_wb_adr_i),
		.userSpace_wb_data_i(userSpace_wb_data_i),
		.userSpace_wb_ack_o(userSpace_wb_ack_o),
		.userSpace_wb_data_o(userSpace_wb_data_o));

	wire userSpaceEnable = userSpace_wb_adr_i[31:28] == USER_SPACE_ADDRESS;
	reg hostConfigLatch = 1'b0;
	wire hostConfigSelect = userSpaceEnable && userSpace_wb_adr_i[27:24] == HOST_PERIPHERAL_ADDRESS;
	wire hostConfigEnable = hostConfigLatch || hostConfigSelect;

	wire caravelHost_wb_ack_o;
	wire caravelHost_wb_stall_o;
	wire caravelHost_wb_error_o;
	wire[31:0] caravelHost_wb_data_o;

	always @(posedge wb_clk_i) begin
		if (wb_rst_i || !userSpace_wb_cyc_i) hostConfigLatch <= 1'b0;
		else if (hostConfigSelect && userSpace_wb_cyc_i) hostConfigLatch <= 1'b1;
	end

	// Caravel wishbone master
	wire caravelEnable = userSpace_wb_cyc_i && userSpaceEnable && !hostConfigEnable;
	assign caravel_wb_cyc_o = caravelEnable;
	assign caravel_wb_stb_o = userSpace_wb_stb_i && caravelEnable;
	assign caravel_wb_we_o = userSpace_wb_we_i && caravelEnable;
	assign caravel_wb_sel_o = caravelEnable ? userSpace_wb_sel_i : 4'b0000;
	assign caravel_wb_data_o = caravelEnable ? userSpace_wb_data_i : ~32'b0;
	assign caravel_wb_adr_o = caravelEnable ? userSpace_wb_adr_i[27:0] : 28'b0;

	always @(*) begin
		if (userSpace_wb_cyc_i) begin
			if (hostConfigEnable) userSpace_wb_ack_o <= caravelHost_wb_ack_o;
			else begin
				if (userSpaceEnable) userSpace_wb_ack_o <= caravel_wb_ack_i || caravel_wb_error_i;
				else userSpace_wb_ack_o <= 1'b1;
			end 
		end else begin
			userSpace_wb_ack_o <= 1'b0;
		end
	end

	//assign userSpace_wb_stall_i = hostConfigEnable ? caravelHost_wb_stall_o : caravel_wb_stall_i;
	//assign userSpace_wb_error_i = hostConfigEnable ? caravelHost_wb_error_o : caravel_wb_error_i;
	assign userSpace_wb_data_o  = hostConfigEnable ? caravelHost_wb_data_o : caravel_wb_data_i;

	// Peripheral bus
	wire peripheralBus_we;
	wire peripheralBus_oe;
	wire peripheralBus_busy;
	wire[23:0] peripheralBus_address;
	wire[3:0] peripheralBus_byteSelect;
	wire[31:0] peripheralBus_dataRead;
	wire[31:0] peripheralBus_dataWrite;
	WBPeripheralBusInterface wbPeripheralBusInterface(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_stb_i(userSpace_wb_stb_i && hostConfigEnable),
		.wb_cyc_i(userSpace_wb_cyc_i && hostConfigEnable),
		.wb_we_i(userSpace_wb_we_i),
		.wb_sel_i(userSpace_wb_sel_i),
		.wb_data_i(userSpace_wb_data_i),
		.wb_adr_i(userSpace_wb_adr_i[23:0]),
		.wb_ack_o(caravelHost_wb_ack_o),
		.wb_stall_o(caravelHost_wb_stall_o),
		.wb_error_o(caravelHost_wb_error_o),
		.wb_data_o(caravelHost_wb_data_o),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(peripheralBus_busy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(peripheralBus_dataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite));

	// Peripheral select
	wire[15:0] localAddress;
	wire peripheralEnable;
	PeripheralSelect #(.ID(4'h0)) select(
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.peripheralEnable(peripheralEnable));

	// UART host
	wire uartOutputRequest_nc;
	wire uartEnable_nc;
	UARTDevice #(.ID(4'h1)) device(
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.peripheralEnable(peripheralEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(peripheralBus_busy),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(peripheralBus_dataRead),
		.requestOutput(uartOutputRequest_nc),
		.uart_en(uartEnable_nc),
		.uart_rx(caravel_uart_rx),
		.uart_tx(caravel_uart_tx));
	
	assign caravel_irq = 3'b0;
	
	assign la_data_out = {
		30'b0,
		probe_out
	};

endmodulemodule WBAddressExtension (
		input wire wb_clk_i,
		input wire wb_rst_i,
		
		// Wishbone Slave port from caravel
		input wire wbs_cyc_i,
		input wire wbs_stb_i,
		input wire wbs_we_i,
		input wire[3:0] wbs_sel_i,
		input wire[31:0] wbs_adr_i,
		input wire[31:0] wbs_data_i,
		output reg wbs_ack_o,
		output reg[31:0] wbs_data_o,

		// Wishbone connection to user space
		output wire userSpace_wb_cyc_i,
		output wire userSpace_wb_stb_i,
		output wire userSpace_wb_we_i,
		output wire[3:0] userSpace_wb_sel_i,
		output wire[31:0] userSpace_wb_adr_i,
		output wire[31:0] userSpace_wb_data_i,
		input wire userSpace_wb_ack_o,
		input wire[31:0] userSpace_wb_data_o
	);
	
	reg[31:0] currentAddress = 32'b0;

	// Connect user space wishbone bus
	wire busAccess = wbs_cyc_i && wbs_adr_i[31:16] == 16'h3000;
	wire userSpaceSelect = busAccess && wbs_adr_i[15];
	wire[14:0] addressOffset = wbs_adr_i[14:0];

	assign userSpace_wb_cyc_i = userSpaceSelect ? wbs_cyc_i : 1'b0;
	assign userSpace_wb_stb_i = userSpaceSelect ? wbs_stb_i : 1'b0;
	assign userSpace_wb_we_i = userSpaceSelect ? wbs_we_i : 1'b0;
	assign userSpace_wb_sel_i = userSpaceSelect ? wbs_sel_i : 4'b0000;
	assign userSpace_wb_adr_i = userSpaceSelect ? { currentAddress[31:15], addressOffset } : 32'b0;
	assign userSpace_wb_data_i = userSpaceSelect ? wbs_data_i : 32'b0;

	// Wishbone interface to allow setting current addres
	localparam STATE_IDLE  		  = 2'h0;
	localparam STATE_WRITE_SINGLE = 2'h1;
	localparam STATE_READ_SINGLE  = 2'h2;
	localparam STATE_FINISH 	  = 2'h3;
	
	reg[1:0] state = STATE_IDLE;
	reg[3:0] currentByteSelect;
	reg[31:0] currentDataIn;

	reg acknowledge = 1'b0;
	reg[31:0] dataRead_buffered = ~32'b0;

	always @(posedge wb_clk_i) begin
		if (wb_rst_i) begin
			state <= STATE_IDLE;
			acknowledge <= 1'b0;
			dataRead_buffered <= ~32'b0;
		end else begin
			case (state)
				STATE_IDLE: begin
					acknowledge <= 1'b0;
					dataRead_buffered <= ~32'b0;

					if (wbs_cyc_i && busAccess && !userSpaceSelect) begin
						if (wbs_stb_i) begin
							if (wbs_we_i) begin
								state <= STATE_WRITE_SINGLE;
							end else begin
								state <= STATE_READ_SINGLE;
							end
						end
					end
				end

				STATE_WRITE_SINGLE: begin
					state <= STATE_FINISH;
					acknowledge <= 1'b1;
					if (wbs_sel_i[0]) currentAddress[7:0]   <= wbs_data_i[7:0];
					if (wbs_sel_i[1]) currentAddress[15:8]  <= wbs_data_i[15:8];
					if (wbs_sel_i[2]) currentAddress[23:16] <= wbs_data_i[23:16];
					if (wbs_sel_i[3]) currentAddress[31:24] <= wbs_data_i[31:24];
				end

				STATE_READ_SINGLE: begin
					state <= STATE_FINISH;
					acknowledge <= 1'b1;
					dataRead_buffered <= currentAddress;
				end

				STATE_FINISH: begin
					state <= STATE_IDLE;
					acknowledge <= 1'b0;
					dataRead_buffered <= ~32'b0;
				end

				default: begin
					state <= STATE_IDLE;
					acknowledge <= 1'b0;
				end				
			endcase
		end
	end

	// Connect wishbone return signals
	always @(*) begin
		if (busAccess) begin
			if (userSpaceSelect) begin
				wbs_ack_o <= userSpace_wb_ack_o;
				wbs_data_o <= userSpace_wb_data_o;
			end else begin
				wbs_ack_o <= acknowledge;
				wbs_data_o <= dataRead_buffered;
			end
		end else begin
			wbs_ack_o <= 1'b0;
			wbs_data_o <= 32'b0;
		end
	end
	
endmodulemodule ExperiarCore (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		input wire wb_clk_i,
		input wire wb_rst_i,

		input wire[7:0] coreIndex,
		input wire[10:0] manufacturerID,
		input wire[15:0] partID,
		input wire[3:0] versionID,

		// JTAG interface
		input wire jtag_tck,
		input wire jtag_tms,
		input wire jtag_tdi,
		output wire jtag_tdo,

		// Interrupts
		input wire[15:0] irq,

		// Wishbone master interface from core
		output wire core_wb_cyc_o,
		output wire core_wb_stb_o,
		output wire core_wb_we_o,
		output wire[3:0] core_wb_sel_o,
		output wire[31:0] core_wb_data_o,
		output wire[27:0] core_wb_adr_o,
		input wire core_wb_ack_i,
		input wire core_wb_stall_i,
		input wire core_wb_error_i,
		input wire[31:0] core_wb_data_i,

		// Wishbone slave interface to sram
		input wire localMemory_wb_cyc_i,
		input wire localMemory_wb_stb_i,
		input wire localMemory_wb_we_i,
		input wire[3:0] localMemory_wb_sel_i,
		input wire[31:0] localMemory_wb_data_i,
		input wire[23:0] localMemory_wb_adr_i,
		output wire localMemory_wb_ack_o,
		output wire localMemory_wb_stall_o,
		output wire localMemory_wb_error_o,
		output wire[31:0] localMemory_wb_data_o,

		// SRAM rw port
		output wire clk0, // Port clock
		output wire[1:0] csb0, // active low chip select
		output wire web0, // active low write control
		output wire[3:0] wmask0, // write mask
		output wire[SRAM_ADDRESS_SIZE-1:0] addr0,
		output wire[31:0] din0,
		input  wire[63:0] dout0,

		// SRAM r port
		output wire clk1,
		output wire[1:0] csb1,
		output wire[SRAM_ADDRESS_SIZE-1:0] addr1,
		input  wire[63:0] dout1,

		// Logic probes
		output wire probe_state,
		output wire[1:0] probe_env,
		output wire[31:0] probe_programCounter,
		output wire[4:0] probe_jtagInstruction
	);
	
	localparam SRAM_ADDRESS_SIZE = 9;

	// Management
	// Shortened form of misa register
	// Modified extensions encounding
	// Origional Bit | New Bit | Character | Description
	// --------------|---------|-----------|------------------------------------------------------
	// 0 			 | 0 	   | A 		   | Atomic extension
	// 1 			 | 1 	   | B 		   | Tentatively reserved for Bit-Manipulation extension
	// 2 			 | 2 	   | C 		   | Compressed extension
	// 3 			 | 3 	   | D 		   | Double-precision floating-point extension
	// 4 			 | 4 	   | E 		   | RV32E base ISA
	// 5 			 | 5 	   | F 		   | Single-precision floating-point extension
	// 6 			 | 6 	   | G 		   | Additional standard extensions present
	// 7 			 | 7 	   | H 		   | Hypervisor extension
	// 8 			 | 8 	   | I 		   | RV32I/64I/128I base ISA
	// 12			 | 9 	   | M 		   | Integer Multiply/Divide extension
	// 13			 | 10 	   | N 		   | User-level interrupts supported
	// 16			 | 11 	   | Q 		   | Quad-precision floating-point extension
	// 18			 | 12 	   | S 		   | Supervisor mode implemented
	// 20			 | 13 	   | U 		   | User mode implemented
	localparam CORE_MXL = 2'h1;
	localparam CORE_EXTENSIONS = 26'b00_0000_0000_0000_0001_0000_0000;
	localparam CORE_EXTENSIONS_SHORT = 14'b00_0001_0000_0000;
	localparam CORE_VERSION = 8'h00;

	// Core
	// Instruction cache interface
	wire[31:0] coreInstructionMemoryAddress;
	wire coreInstructionMemoryEnable;
	wire[31:0] coreInstructionMemoryDataRead;
	wire coreInstructionMemoryBusy;
	wire coreInstructionMemoryAccessFault = |(coreInstructionMemoryAddress[1:0]);
	wire coreInstructionAddressBreakpoint;

	// Data cache interface
	wire[31:0] coreDataMemoryAddress;
	wire[3:0] coreDataMemoryByteSelect;
	wire coreDataMemoryEnable;
	wire coreDataMemoryWriteEnable;
	wire[31:0] coreDataMemoryDataWrite;
	wire[31:0] coreDataMemoryDataRead;
	wire coreDataMemoryBusy;
	wire coreDataMemoryAccessFault = |(coreDataMemoryAddress[1:0]);
	wire coreDataAddressBreakpoint;

	// Memory interface from core to local memory
	wire coreLocalMemoryEnable;
	wire coreLocalMemoryWriteEnable;
	wire[23:0] coreLocalMemoryAddress;
	wire[3:0] coreLocalMemoryByteSelect;
	wire[31:0] coreLocalMemoryDataWrite;
	wire[31:0] coreLocalMemoryDataRead;
	wire coreLocalMemoryBusy;

	// Memory interface from core to wb
	wire coreWBEnable;
	wire coreWBWriteEnable;
	wire[27:0] coreWBAddress;
	wire[3:0] coreWBByteSelect;
	wire[31:0] coreWBDataWrite;
	wire[31:0] coreWBDataRead;
	wire coreWBBusy;

	// Memory interface from wb to local memory
	wire wbLocalMemoryEnable;
	wire wbLocalMemoryWriteEnable;
	wire[23:0] wbLocalMemoryAddress;
	wire[3:0] wbLocalMemoryByteSelect;
	wire[31:0] wbLocalMemoryDataWrite;
	wire[31:0] wbLocalMemoryDataRead;
	wire wbLocalMemoryBusy;

	// Core management
	wire management_run;
	wire management_interruptEnable;
	wire management_writeEnable;
	wire[3:0] management_byteSelect;
	wire[15:0] management_address;
	wire[31:0] management_writeData;
	wire[31:0] management_readData;

	wire jtag_management_enable;
	wire jtag_management_writeEnable;
	wire[3:0] jtag_management_byteSelect;
	wire[19:0] jtag_management_address;
	wire[31:0] jtag_management_writeData;
	wire[31:0] jtag_management_readData;

	wire wb_management_enable;
	wire wb_management_writeEnable;
	wire[3:0] wb_management_byteSelect;
	wire[19:0] wb_management_address;
	wire[31:0] wb_management_writeData;
	wire[31:0] wb_management_readData;
	wire wb_management_busy;

	JTAG jtag(
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.coreID({ coreIndex, CORE_VERSION, CORE_MXL, CORE_EXTENSIONS_SHORT }),
		.manufacturerID(manufacturerID),
		.partID(partID),
		.versionID(versionID),
		.jtag_tck(jtag_tck),
		.jtag_tms(jtag_tms),
		.jtag_tdi(jtag_tdi),
		.jtag_tdo(jtag_tdo),
		.management_enable(jtag_management_enable),
		.management_writeEnable(jtag_management_writeEnable),
		.management_byteSelect(jtag_management_byteSelect),
		.management_address(jtag_management_address),
		.management_writeData(jtag_management_writeData),
		.management_readData(jtag_management_readData),
		.probe_jtagInstruction(probe_jtagInstruction));

	CoreManagement coreManagement(
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.management_run(management_run),
		.management_interruptEnable(management_interruptEnable),
		.management_writeEnable(management_writeEnable),
		.management_byteSelect(management_byteSelect),
		.management_address(management_address),
		.management_writeData(management_writeData),
		.management_readData(management_readData),
		.isInstructionAddressBreakpoint(coreInstructionAddressBreakpoint),
		.isDataAddressBreakpoint(coreDataAddressBreakpoint),
		.coreInstructionAddress(coreInstructionMemoryAddress),
		.coreDataAddress(coreDataMemoryAddress),
		.jtag_management_enable(jtag_management_enable),
		.jtag_management_writeEnable(jtag_management_writeEnable),
		.jtag_management_byteSelect(jtag_management_byteSelect),
		.jtag_management_address(jtag_management_address),
		.jtag_management_writeData(jtag_management_writeData),
		.jtag_management_readData(jtag_management_readData),
		.wb_management_enable(wb_management_enable),
		.wb_management_writeEnable(wb_management_writeEnable),
		.wb_management_byteSelect(wb_management_byteSelect),
		.wb_management_address(wb_management_address),
		.wb_management_writeData(wb_management_writeData),
		.wb_management_readData(wb_management_readData),
		.wb_management_busy(wb_management_busy));

	// Core
	RV32ICore core(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.instruction_memoryAddress(coreInstructionMemoryAddress),
		.instruction_memoryEnable(coreInstructionMemoryEnable),
		.instruction_memoryDataRead(coreInstructionMemoryDataRead),
		.instruction_memoryBusy(coreInstructionMemoryBusy),
		.instruction_memoryAccessFault(coreInstructionMemoryAccessFault),
		.instruction_memoryAddressBreakpoint(coreInstructionAddressBreakpoint),
		.data_memoryAddress(coreDataMemoryAddress),
		.data_memoryByteSelect(coreDataMemoryByteSelect),
		.data_memoryEnable(coreDataMemoryEnable),
		.data_memoryWriteEnable(coreDataMemoryWriteEnable),
		.data_memoryDataWrite(coreDataMemoryDataWrite),
		.data_memoryDataRead(coreDataMemoryDataRead),
		.data_memoryBusy(coreDataMemoryBusy),
		.data_memoryAccessFault(coreDataMemoryAccessFault),
		.data_memoryAddressBreakpoint(coreDataAddressBreakpoint),
		.management_run(management_run),
		.management_interruptEnable(management_interruptEnable),
		.management_writeEnable(management_writeEnable),
		.management_byteSelect(management_byteSelect),
		.management_address(management_address),
		.management_writeData(management_writeData),
		.management_readData(management_readData),
		.coreIndex(coreIndex),
		.manufacturerID(manufacturerID),
		.partID(partID),
		.versionID(versionID),
		.extensions(CORE_EXTENSIONS),
		.userInterrupts(irq),
		.probe_state(probe_state),
		.probe_env(probe_env),
		.probe_programCounter(probe_programCounter));

	MemoryController memoryController(
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.coreInstructionAddress(coreInstructionMemoryAddress),
		.coreInstructionEnable(coreInstructionMemoryEnable),
		.coreInstructionDataRead(coreInstructionMemoryDataRead),
		.coreInstructionBusy(coreInstructionMemoryBusy),
		.coreDataAddress(coreDataMemoryAddress),
		.coreDataByteSelect(coreDataMemoryByteSelect),
		.coreDataEnable(coreDataMemoryEnable),
		.coreDataWriteEnable(coreDataMemoryWriteEnable),
		.coreDataDataWrite(coreDataMemoryDataWrite),
		.coreDataDataRead(coreDataMemoryDataRead),
		.coreDataBusy(coreDataMemoryBusy),
		.localMemoryAddress(coreLocalMemoryAddress),
		.localMemoryByteSelect(coreLocalMemoryByteSelect),
		.localMemoryWriteEnable(coreLocalMemoryWriteEnable),
		.localMemoryEnable(coreLocalMemoryEnable),
		.localMemoryDataWrite(coreLocalMemoryDataWrite),
		.localMemoryDataRead(coreLocalMemoryDataRead),
		.localMemoryBusy(coreLocalMemoryBusy),
		.wbAddress(coreWBAddress),
		.wbByteSelect(coreWBByteSelect),
		.wbEnable(coreWBEnable),
		.wbWriteEnable(coreWBWriteEnable),
		.wbDataWrite(coreWBDataWrite),
		.wbDataRead(coreWBDataRead),
		.wbBusy(coreWBBusy));

	LocalMemoryInterface #(.SRAM_ADDRESS_SIZE(SRAM_ADDRESS_SIZE)) localMemoryInterface (
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.coreAddress(coreLocalMemoryAddress),
		.coreByteSelect(coreLocalMemoryByteSelect),
		.coreEnable(coreLocalMemoryEnable),
		.coreWriteEnable(coreLocalMemoryWriteEnable),
		.coreDataWrite(coreLocalMemoryDataWrite),
		.coreDataRead(coreLocalMemoryDataRead),
		.coreBusy(coreLocalMemoryBusy),
		.wbAddress(wbLocalMemoryAddress),
		.wbByteSelect(wbLocalMemoryByteSelect),
		.wbEnable(wbLocalMemoryEnable),
		.wbWriteEnable(wbLocalMemoryWriteEnable),
		.wbDataWrite(wbLocalMemoryDataWrite),
		.wbDataRead(wbLocalMemoryDataRead),
		.wbBusy(wbLocalMemoryBusy),
		.clk0(clk0),
		.csb0(csb0),
		.web0(web0),
		.wmask0(wmask0),
		.addr0(addr0),
		.din0(din0),
		.dout0(dout0),
		.clk1(clk1),
		.csb1(csb1),
		.addr1(addr1),
		.dout1(dout1));

	Core_WBInterface coreWBInterface(
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_cyc_o(core_wb_cyc_o),
		.wb_stb_o(core_wb_stb_o),
		.wb_we_o(core_wb_we_o),
		.wb_sel_o(core_wb_sel_o),
		.wb_data_o(core_wb_data_o),
		.wb_adr_o(core_wb_adr_o),
		.wb_ack_i(core_wb_ack_i),
		.wb_stall_i(core_wb_stall_i),
		.wb_error_i(core_wb_error_i),
		.wb_data_i(core_wb_data_i),
		.wbAddress(coreWBAddress),
		.wbByteSelect(coreWBByteSelect),
		.wbEnable(coreWBEnable),
		.wbWriteEnable(coreWBWriteEnable),
		.wbDataWrite(coreWBDataWrite),
		.wbDataRead(coreWBDataRead),
		.wbBusy(coreWBBusy));

	WB_SRAMInterface wbSRAMInterface(
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_cyc_i(localMemory_wb_cyc_i),
		.wb_stb_i(localMemory_wb_stb_i),
		.wb_we_i(localMemory_wb_we_i),
		.wb_sel_i(localMemory_wb_sel_i),
		.wb_data_i(localMemory_wb_data_i),
		.wb_adr_i(localMemory_wb_adr_i),
		.wb_ack_o(localMemory_wb_ack_o),
		.wb_stall_o(localMemory_wb_stall_o),
		.wb_error_o(localMemory_wb_error_o),
		.wb_data_o(localMemory_wb_data_o),
		.localMemoryAddress(wbLocalMemoryAddress),
		.localMemoryByteSelect(wbLocalMemoryByteSelect),
		.localMemoryEnable(wbLocalMemoryEnable),
		.localMemoryWriteEnable(wbLocalMemoryWriteEnable),
		.localMemoryDataWrite(wbLocalMemoryDataWrite),
		.localMemoryDataRead(wbLocalMemoryDataRead),
		.localMemoryBusy(wbLocalMemoryBusy),
		.management_enable(wb_management_enable),
		.management_writeEnable(wb_management_writeEnable),
		.management_byteSelect(wb_management_byteSelect),
		.management_address(wb_management_address),
		.management_writeData(wb_management_writeData),
		.management_readData(wb_management_readData),
		.management_busy(wb_management_busy));

endmodulemodule CoreManagement (
		input wire clk,
		input wire rst,

		// Interface to core
		output wire management_run,
		output wire management_interruptEnable,
		output wire management_writeEnable,
		output wire[3:0] management_byteSelect,
		output wire[15:0] management_address,
		output wire[31:0] management_writeData,
		input wire[31:0] management_readData,

		// Address breakpoint
		output wire isInstructionAddressBreakpoint,
		output wire isDataAddressBreakpoint,
		input wire[31:0] coreInstructionAddress,
		input wire[31:0] coreDataAddress,

		// Interface from jtag
		input wire jtag_management_enable,
		input wire jtag_management_writeEnable,
		input wire[3:0] jtag_management_byteSelect,
		input wire[19:0] jtag_management_address,
		input wire[31:0] jtag_management_writeData,
		output wire[31:0] jtag_management_readData,

		// Interface from wishbone
		input wire wb_management_enable,
		input wire wb_management_writeEnable,
		input wire[3:0] wb_management_byteSelect,
		input wire[19:0] wb_management_address,
		input wire[31:0] wb_management_writeData,
		output wire[31:0] wb_management_readData,
		output wire wb_management_busy
	);

	// TODO instruction breakpoints
	assign isInstructionAddressBreakpoint = 0;
	assign isDataAddressBreakpoint = 0;
	//assign isInstructionAddressBreakpoint = coreInstructionAddress == instructionBreakpointAddress;
	//assign isDataAddressBreakpoint = coreDataAddress == dataBreakpointAddress;

	// Master select
	wire jtagSelect = jtag_management_enable;
	wire wbRequest = wb_management_enable;
	wire wbSelect = wbRequest && !jtagSelect;

	wire peripheralBus_we = jtag_management_writeEnable || (!jtagSelect && wb_management_writeEnable);
	wire peripheralBus_oe = (jtag_management_enable && !jtag_management_writeEnable)  || (!jtagSelect && wb_management_enable && !wb_management_writeEnable);
	wire[19:0] peripheralBus_address = jtagSelect ? jtag_management_address : 
								   	   wbSelect   ? wb_management_address   : 20'b0;
	wire[3:0] peripheralBus_byteSelect = jtagSelect ? jtag_management_byteSelect : 
								   	     wbSelect   ? wb_management_byteSelect   : 4'h0;
	wire[31:0] peripheralBus_dataWrite = jtag_management_writeEnable ? jtag_management_writeData :
									 	 wb_management_writeEnable   ? wb_management_writeData   : 32'b0;

	wire[31:0] peripheralBus_dataRead;
	assign jtag_management_readData = peripheralBus_dataRead;
	assign wb_management_readData = peripheralBus_dataRead;
	assign wb_management_busy = jtagSelect && wbRequest;

	wire registerEnable = peripheralBus_address[19:12] == 8'h00;
	wire coreEnable = peripheralBus_address[19:16] == 4'h1 && !management_run;

	// Registers
	// Control register: Default 0x0
	// b00: run
	// b01: unused
	// b02: interruptEnable
	wire[2:0] control;
	wire[31:0] controlOutputData;
	wire controlOutputRequest;
	ConfigurationRegister #(.WIDTH(3), .ADDRESS(12'h000), .DEFAULT(3'b0)) controlRegister(
		.clk(clk),
		.rst(rst),
		.enable(registerEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(peripheralBus_address[11:0]),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(controlOutputData),
		.requestOutput(controlOutputRequest),
		.currentValue(control));

	// Core
	assign management_run = control[0];
	assign management_interruptEnable = control[2];
	assign management_writeEnable = coreEnable && peripheralBus_we;
	assign management_byteSelect = peripheralBus_byteSelect;
	assign management_address = peripheralBus_address[15:0];
	assign management_writeData = peripheralBus_dataWrite;

	assign peripheralBus_dataRead = coreEnable 			 ? management_readData :
									controlOutputRequest ? controlOutputData   : ~32'b0;
	
endmodulemodule RV32ICore(

	inout vccd1,	// User area 1 1.8V supply
	inout vssd1,	// User area 1 digital ground


		input wire clk,
		input wire rst,

		// Instruction cache interface
		output wire[31:0] instruction_memoryAddress,
		output wire instruction_memoryEnable,
		input wire[31:0] instruction_memoryDataRead,
		input wire instruction_memoryBusy,
		input wire instruction_memoryAccessFault,
		input wire instruction_memoryAddressBreakpoint,

		// Data cache interface
		output wire[31:0] data_memoryAddress,
		output wire[3:0] data_memoryByteSelect,
		output wire data_memoryEnable,
		output wire data_memoryWriteEnable,
		output wire[31:0] data_memoryDataWrite,
		input wire[31:0] data_memoryDataRead,
		input wire data_memoryBusy,
		input wire data_memoryAccessFault,
		input wire data_memoryAddressBreakpoint,

		// Management interface
		input wire management_run,
		input wire management_interruptEnable,
		input wire management_writeEnable,
		input wire[3:0] management_byteSelect,
		input wire[15:0] management_address,
		input wire[31:0] management_writeData,
		output wire[31:0] management_readData,

		// System info
		input wire[7:0] coreIndex,
		input wire[10:0] manufacturerID,
		input wire[15:0] partID,
		input wire[3:0] versionID,
		input wire[25:0] extensions,

		// Traps
		input wire[15:0] userInterrupts,

		// Logic probes
		output wire probe_state,
		output wire[1:0] probe_env,
		output wire[31:0] probe_programCounter
    );

	localparam STATE_HALT 	 	= 1'b0;
	localparam STATE_EXECUTE 	= 1'b1;

	//localparam STATE_HALT 	 	= 2'b00;
	//localparam STATE_FETCH   	= 2'b10;
	//localparam STATE_EXECUTE 	= 2'b11;

	// System registers
	reg state = STATE_HALT;
	reg[31:0] fetchProgramCounter = 32'b0;
	reg[31:0] executeProgramCounter = 32'b0;
	reg[31:0] registers [0:31];

	// Management control
	localparam MANAGMENT_ADDRESS_SYSTEM	   = 2'b00;
	localparam MANAGMENT_ADDRESS_REGISTERS = 2'b01;
	localparam MANAGMENT_ADDRESS_CSR 	   = 2'b10;

	wire management_selectProgramCounter      = (management_address[15:14] == MANAGMENT_ADDRESS_SYSTEM) && (management_address[13:4] == 10'h000);
	wire management_selectInstructionRegister = (management_address[15:14] == MANAGMENT_ADDRESS_SYSTEM) && (management_address[13:4] == 10'h001);
	wire management_selectClearError		  = (management_address[15:14] == MANAGMENT_ADDRESS_SYSTEM) && (management_address[13:4] == 10'h002);
	wire management_selectRegister            = (management_address[15:14] == MANAGMENT_ADDRESS_REGISTERS) && (management_address[13:7] == 7'h00);
	wire management_selectCSR 				  = management_address[15:14] == MANAGMENT_ADDRESS_CSR;

	wire management_writeValid = !management_run && management_writeEnable;
	wire management_writeProgramCounter = management_writeValid && management_selectProgramCounter;
	wire management_writeProgramCounter_set = management_writeProgramCounter && (management_address[3:0] == 4'h0);
	wire management_writeProgramCounter_jump = management_writeProgramCounter && (management_address[3:0] == 4'h4);
	wire management_writeProgramCounter_step = management_writeProgramCounter && (management_address[3:0] == 4'h8);
	wire management_writeClearError = management_writeValid && management_selectClearError;
	wire management_writeRegister = management_writeValid && management_selectRegister;
	wire management_writeCSR = management_writeValid && management_selectCSR;

	wire management_readValid = !management_run && !management_writeEnable;
	wire management_readProgramCounter = management_readValid && management_selectProgramCounter;
	wire management_readInstructionRegister = management_readValid && management_selectInstructionRegister;
	wire management_readRegister = management_readValid && management_selectRegister;
	wire management_readCSR = management_readValid && management_selectCSR;

	wire pipeActive;
	reg stepProgramCounter;

	// Make sure to flush the pipe after a step
	reg management_pipeStartup = 1'b0;
	always @(posedge clk) begin
		if (rst) begin
			management_pipeStartup <= 1'b0;
		end else begin
			if ((management_run || management_writeProgramCounter_step) && !management_pipeStartup) management_pipeStartup <= 1'b1;
			else if (stepProgramCounter) management_pipeStartup <= 1'b0;
		end
	end

	wire management_allowInstruction = management_run || management_writeProgramCounter_step || management_pipeStartup;

	wire[4:0] management_registerIndex = management_address[6:2];
	wire[11:0] management_csrIndex = management_address[13:2];

	reg[31:0] management_dataOut;

	wire[31:0] csrReadData;

	always @(*) begin
		case (1'b1)
			management_readProgramCounter: management_dataOut <= fetchProgramCounter;
			management_readInstructionRegister : management_dataOut <= pipe1_currentInstruction;
			management_readRegister: management_dataOut <= !management_registerIndex ? registers[management_registerIndex] : 32'b0;
			management_readCSR: management_dataOut <= csrReadData;
			default: management_dataOut <= ~32'b0;
		endcase
	end

	assign management_readData = {
		management_byteSelect[3] ? management_dataOut[31:24] : 8'h00,
		management_byteSelect[2] ? management_dataOut[23:16] : 8'h00,
		management_byteSelect[1] ? management_dataOut[15:8]  : 8'h00,
		management_byteSelect[0] ? management_dataOut[7:0]   : 8'h00
	};

	wire[31:0] trapVector;
	wire[31:0] trapReturnVector;
	wire inTrap;

	// ----------Pipe----------
	wire pipe1_shouldStall;
	wire pipe2_shouldStall;
	wire shouldStore;
	wire shouldLoad;

	reg cancelStall;

	wire loadStoreBusy = shouldStore || shouldLoad ? data_memoryBusy : 1'b0;
	wire stepBlocked = (instruction_memoryEnable && instruction_memoryBusy) || loadStoreBusy;// || !management_allowInstruction
	wire stepPipe = state == STATE_EXECUTE && !stepBlocked;
	wire progressPipe = pipeActive || management_allowInstruction;
	wire stallPipe = !management_allowInstruction || pipe1_shouldStall || pipe2_shouldStall;
	wire stallIncrementProgramCounter = !management_allowInstruction || pipe1_shouldStall;

	// 0: Request instruction
	wire pipe0_stall;
	wire pipe0_active;
	wire[31:0] pipe0_currentInstruction;
	wire[31:0] pipe0_programCounter;
	wire pipe0_addressMisaligned;
	wire[31:0] pipe0_instructionFetchAddress;
	wire pipe0_instructionFetchEnable;
	PipeFetch pipe0_fetch (
		.clk(clk),
		.rst(rst),
		.stepPipe(stepPipe),
		.pipeStall(stallPipe),
		.currentPipeStall(pipe0_stall),
		.active(pipe0_active),
		.currentInstruction(instruction_memoryDataRead),
		.lastInstruction(pipe0_currentInstruction),
		.programCounter(fetchProgramCounter),
		.lastProgramCounter(pipe0_programCounter),
		.addressMisaligned(pipe0_addressMisaligned),
		.fetchAddress(pipe0_instructionFetchAddress),
		.fetchEnable(pipe0_instructionFetchEnable));

	// 1: Request data/Write data/ALU operation
	reg[31:0] pipe1_resultRegister;
	reg[31:0] pipe1_csrData;

	wire pipe1_stall;
	wire pipe1_active;
	wire pipe1_invalidInstruction;
	wire[31:0] pipe1_currentInstruction;
	wire[11:0] pipe1_csrReadAddress;
	wire pipe1_csrReadEnable;

	wire[4:0] pipe1_rs1Address;
	wire[4:0] pipe1_rs2Address;
	reg[31:0] pipe1_rs1Data;
	reg[31:0] pipe1_rs2Data;
	wire pipe1_operationResultStoreEnable;
	wire[31:0] pipe1_operationResult;
	wire pipe1_isJump;
	wire pipe1_isFence;
	wire pipe1_jumpEnable;
	wire pipe1_failedBranch;
	wire[31:0] pipe1_nextProgramCounter;
	wire pipe1_jumpMissaligned;
	wire pipe1_addressMisaligned_load;
	wire pipe1_addressMisaligned_store;
	wire pipe1_memoryEnable;
	wire pipe1_memoryWriteEnable;
	wire[3:0] pipe1_memoryByteSelect;
	wire[31:0] pipe1_memoryAddress;
	wire[31:0] pipe1_memoryWriteData;
	wire[31:0] pipe1_fullMemoryAddress;
	wire pipe1_isECALL;
	wire pipe1_isEBREAK;
	wire pipe1_isRET;
	PipeOperation pipe1_operation (
		.clk(clk),
		.rst(rst),
		.stepPipe(stepPipe),
		.pipeStall(pipe0_stall && !cancelStall),
		.currentPipeStall(pipe1_stall),
		.active(pipe1_active),
		.currentInstruction(pipe0_currentInstruction),
		.lastInstruction(pipe1_currentInstruction),
		.invalidInstruction(pipe1_invalidInstruction),
		.csrReadAddress(pipe1_csrReadAddress),
		.csrReadData(csrReadData),
		.csrReadEnable(pipe1_csrReadEnable),
		.programCounter(executeProgramCounter),
		.rs1Address(pipe1_rs1Address),
		.rs1Data(pipe1_rs1Data),
		.rs2Address(pipe1_rs2Address),
		.rs2Data(pipe1_rs2Data),
		.operationResultStoreEnable(pipe1_operationResultStoreEnable),
		.operationResult(pipe1_operationResult),
		.isJump(pipe1_isJump),
		.isFence(pipe1_isFence),
		.jumpEnable(pipe1_jumpEnable),
		.failedBranch(pipe1_failedBranch),
		.nextProgramCounter(pipe1_nextProgramCounter),
		.jumpMissaligned(pipe1_jumpMissaligned),
		.addressMisaligned_load(pipe1_addressMisaligned_load),
		.addressMisaligned_store(pipe1_addressMisaligned_store),
		.memoryEnable(pipe1_memoryEnable),
		.memoryWriteEnable(pipe1_memoryWriteEnable),
		.memoryByteSelect(pipe1_memoryByteSelect),
		.memoryAddress(pipe1_memoryAddress),
		.memoryWriteData(pipe1_memoryWriteData),
		.fullMemoryAddress(pipe1_fullMemoryAddress),
		.isECALL(pipe1_isECALL),
		.isEBREAK(pipe1_isEBREAK),
		.isRET(pipe1_isRET));

	assign pipe1_shouldStall = pipe1_isJump || pipe1_isFence || pipe1_isRET;

	always @(posedge clk) begin
		if (rst) begin
			pipe1_resultRegister <= 32'b0;
			pipe1_csrData <= 32'b0;
			cancelStall <= 1'b0;
		end else begin
			if (state == STATE_EXECUTE) begin
				if (pipe1_operationResultStoreEnable) pipe1_resultRegister <= pipe1_operationResult;
				if (pipe1_csrReadEnable) pipe1_csrData <= csrReadData;
				cancelStall <= pipe1_failedBranch;
			end
		end
	end

	// 3: Store data
	wire pipe2_stall;
	wire pipe2_active;
	wire pipe2_invalidInstruction;
	wire[31:0] pipe2_currentInstruction;
	wire pipe2_expectingLoad;
	wire[4:0] pipe2_rdAddress;
	wire[31:0] pipe2_registerWriteData;
	wire pipe2_registerWriteEnable;
	wire[11:0] pipe2_csrWriteAddress;
	wire[31:0] pipe2_csrWriteData;
	wire pipe2_csrWriteEnable;
	wire pipe2_isJump;
	wire pipe2_isFence;
	wire pipe2_isRET;
	PipeStore pipe2_store (
		.clk(clk),
		.rst(rst),
		.stepPipe(stepPipe),
		.pipeStall(pipe1_stall),
		.currentPipeStall(pipe2_stall),
		.active(pipe2_active),
		.currentInstruction(pipe1_currentInstruction),
		.lastInstruction(pipe2_currentInstruction),
		.invalidInstruction(pipe2_invalidInstruction),
		.expectingLoad(pipe2_expectingLoad),
		.memoryDataRead(data_memoryDataRead),
		.aluResultData(pipe1_resultRegister),
		.csrData(pipe1_csrData),
		.registerWriteAddress(pipe2_rdAddress),
		.registerWriteData(pipe2_registerWriteData),
		.registerWriteEnable(pipe2_registerWriteEnable),
		.csrWriteAddress(pipe2_csrWriteAddress),
		.csrWriteData(pipe2_csrWriteData),
		.csrWriteEnable(pipe2_csrWriteEnable),
		.isJump(pipe2_isJump),
		.isFence(pipe2_isFence),
		.isRET(pipe2_isRET));

	assign pipe2_shouldStall = pipe2_isJump || pipe2_isFence || pipe2_isRET;
	assign pipeActive = pipe0_active || pipe1_active || pipe2_active;

	// Integer restister control
	// Check if pipe1 needs the value being written by pipe2
	always @(*) begin
		if (pipe2_registerWriteEnable && pipe2_rdAddress == pipe1_rs1Address) begin
			pipe1_rs1Data <= |pipe1_rs1Address ? pipe2_registerWriteData : 32'b0;
		end else begin
			pipe1_rs1Data <= |pipe1_rs1Address ? registers[pipe1_rs1Address] : 32'b0;
		end

		if (pipe2_registerWriteEnable && pipe2_rdAddress == pipe1_rs2Address) begin
			pipe1_rs2Data <= |pipe1_rs2Address ? pipe2_registerWriteData : 32'b0;
		end else begin
			pipe1_rs2Data <= |pipe1_rs2Address ? registers[pipe1_rs2Address] : 32'b0;
		end
	end

	always @(posedge clk) begin
		if (rst) begin
		end else begin
			if (state == STATE_EXECUTE) begin
				if (pipe2_registerWriteEnable && |pipe2_rdAddress) registers[pipe2_rdAddress] <= pipe2_registerWriteData;
			end
		end
	end

	assign shouldStore = pipe1_memoryEnable && pipe1_memoryWriteEnable;
	assign shouldLoad = (pipe1_memoryEnable && !pipe1_memoryWriteEnable) || pipe2_expectingLoad;

	reg[31:0] nextFetchProgramCounter;

	always @(*) begin
		if (rst) begin
			nextFetchProgramCounter = 32'b0;
			stepProgramCounter = 1'b0;
		end else begin
			nextFetchProgramCounter = fetchProgramCounter;
			stepProgramCounter = 1'b0;

			case (state)
				STATE_EXECUTE: begin
					if (stepPipe) begin
						if (inTrap) begin
							nextFetchProgramCounter = trapVector;
							stepProgramCounter = 1'b1;
						end	else if (pipe1_isRET) begin
							nextFetchProgramCounter = trapReturnVector;
							stepProgramCounter = 1'b1;
						end else if (pipe1_jumpEnable) begin
							nextFetchProgramCounter = pipe1_nextProgramCounter;
							stepProgramCounter = 1'b1;
						end else if (!stallPipe) begin
							nextFetchProgramCounter = fetchProgramCounter + 4;
							stepProgramCounter = 1'b1;
						end
					end
				end
			endcase
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			state <= STATE_HALT;
			fetchProgramCounter <= 32'b0;
			executeProgramCounter <= 32'b0;
		end else begin
			case (state)
				STATE_HALT: begin
					if (progressPipe) begin
						state <= STATE_EXECUTE;
					end else begin
						if (management_writeProgramCounter_set) fetchProgramCounter <= management_writeData;
						else if (management_writeProgramCounter_jump) fetchProgramCounter <= executeProgramCounter + management_writeData;
					end
				end

				STATE_EXECUTE: begin
					if (stepPipe) begin
						if (!progressPipe) state <= STATE_HALT;
						if (stepProgramCounter) fetchProgramCounter <= nextFetchProgramCounter;
						executeProgramCounter <= pipe0_programCounter;
					end
				end

				default: state <= STATE_HALT;
			endcase
		end
	end

	// Memory control
	assign instruction_memoryAddress = pipe0_instructionFetchAddress;
	assign instruction_memoryEnable = pipe0_instructionFetchEnable;

	assign data_memoryAddress = pipe1_memoryAddress;
	assign data_memoryByteSelect = pipe1_memoryByteSelect;
	assign data_memoryEnable = pipe1_memoryEnable;
	assign data_memoryWriteEnable = pipe1_memoryWriteEnable;
	assign data_memoryDataWrite = pipe1_memoryWriteData;

	// System commands 
	wire eCall = pipe1_isECALL && (state == STATE_EXECUTE);
	wire eBreak = pipe1_isEBREAK && (state == STATE_EXECUTE);
	wire trapReturn = pipe1_isRET && (state == STATE_EXECUTE);

	wire isMachineTimerInterrupt = 1'b0;
	wire isMachineExternalInterrupt = 1'b0;
	wire isMachineSoftwareInterrupt = 1'b0;

	// CSRs
	// CSR interface
	wire csrWriteEnable = management_writeCSR || (management_run && pipe2_csrWriteEnable && (state == STATE_EXECUTE));
	wire csrReadEnable = management_readCSR || (management_run && pipe1_csrReadEnable && (state == STATE_EXECUTE));
	wire[11:0] csrWriteAddress = !management_run ? management_csrIndex : pipe2_csrWriteAddress;
	wire[11:0] csrReadAddress = !management_run ? management_csrIndex : pipe1_csrReadAddress;
	wire[31:0] csrWriteData = !management_run ? management_writeData : pipe2_csrWriteData;
	
	wire instructionCompleted = !pipe2_stall;
	CSR csr(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(csrReadData),
		.coreIndex(coreIndex),
		.manufacturerID(manufacturerID),
		.partID(partID),
		.versionID(versionID),
		.extensions(extensions),
		.instructionCompleted(instructionCompleted),
		.programCounter(executeProgramCounter),
		.currentInstruction(pipe1_currentInstruction),
		.instruction_memoryAddress(instruction_memoryAddress),
		.data_memoryAddress(pipe1_fullMemoryAddress),
		.isMachineTimerInterrupt(isMachineTimerInterrupt),
		.isMachineExternalInterrupt(isMachineExternalInterrupt),
		.isMachineSoftwareInterrupt(isMachineSoftwareInterrupt),
		.isFetchAddressMisaligned(pipe0_addressMisaligned),
		.isDataAddressMisaligned_load(pipe1_addressMisaligned_load),
		.isDataAddressMisaligned_store(pipe1_addressMisaligned_store),
		.isJumpMissaligned(pipe1_jumpMissaligned),
		.isFetchAccessFault(instruction_memoryAccessFault),
		.isDataAccessFault_load(data_memoryAccessFault && data_memoryEnable && !data_memoryWriteEnable),
		.isDataAccessFault_store(data_memoryAccessFault && data_memoryEnable && data_memoryWriteEnable),
		.isInvalidInstruction(pipe1_invalidInstruction),
		.isEBREAK(eBreak),
		.isECALL(eCall),
		.isFetchAddressBreakpoint(instruction_memoryAddressBreakpoint),
		.isDataAddressBreakpoint(data_memoryAddressBreakpoint),
		.userInterrupts(management_interruptEnable ? userInterrupts : 16'b0),
		.trapReturn(trapReturn),
		.inTrap(inTrap),
		.trapVector(trapVector),
		.trapReturnVector(trapReturnVector));

	// Debug
	assign probe_state = state;
	assign probe_env = { eCall, eBreak };
	assign probe_programCounter = executeProgramCounter;

endmodule
module PipeFetch #(
	 	parameter PROGRAM_COUNTER_RESET = 32'b0
	)(
		input wire clk,
		input wire rst,

		// Pipe control
		input wire stepPipe,
		input wire pipeStall,
		output reg currentPipeStall,
		output wire active,
		input wire[31:0] currentInstruction,
		output reg[31:0] lastInstruction,

		// Control
		input wire[31:0] programCounter,
		output reg[31:0] lastProgramCounter,
		output wire addressMisaligned,		

		// Memory access
		output wire[31:0] fetchAddress,
		output wire fetchEnable
	);

	// Pipe control
	always @(posedge clk) begin
		if (rst) begin
			currentPipeStall <= 1'b1;
			lastInstruction <= 32'b0;
		end else begin
			if (stepPipe) begin
				currentPipeStall <= pipeStall;
				if (!pipeStall) lastInstruction <= currentInstruction;
			end
		end
	end

	assign active = !pipeStall;

	always @(posedge clk) begin
		if (rst) lastProgramCounter <= 32'b0;
		else lastProgramCounter <= programCounter;
	end

	assign addressMisaligned = |programCounter[1:0];

	assign fetchAddress = programCounter;
	assign fetchEnable = !pipeStall;//stepPipe;

endmodulemodule PipeOperation (
		input wire clk,
		input wire rst,

		// Pipe control
		input wire stepPipe,
		input wire pipeStall,
		output wire currentPipeStall,
		output wire active,
		input wire[31:0] currentInstruction,
		output wire[31:0] lastInstruction,
		output wire invalidInstruction,

		// CSR read control
		output wire[11:0] csrReadAddress,
		input wire[31:0] csrReadData,
		output wire csrReadEnable,

		// Operation inputs
		input wire[31:0] programCounter,
		output wire[4:0] rs1Address,
		input wire[31:0] rs1Data,
		output wire[4:0] rs2Address,
		input wire[31:0] rs2Data,

		// Operation outputs
		output wire operationResultStoreEnable,
		output wire[31:0] operationResult,
		output wire isJump,
		output wire isFence,
		output wire jumpEnable,
		output wire failedBranch,
		output wire[31:0] nextProgramCounter,
		output wire jumpMissaligned,
		output wire addressMisaligned_load,
		output wire addressMisaligned_store,

		// Load/Store control
		output wire memoryEnable,
		output wire memoryWriteEnable,
		output wire[3:0] memoryByteSelect,
		output wire[31:0] memoryAddress,
		output wire[31:0] memoryWriteData,
		output wire[31:0] fullMemoryAddress,

		// System operations
		output wire isECALL,
		output wire isEBREAK,
		output wire isRET
	);

	// Pipe control
	PipeStage pipeStage(
		.clk(clk),
		.rst(rst),
		.stepPipe(stepPipe),
		.pipeStall(pipeStall),
		.currentPipeStall(currentPipeStall),
		.active(active),
		.currentInstruction(currentInstruction),
		.lastInstruction(lastInstruction));

	// Instruction decode
	wire[6:0] opcode;
	wire[4:0] rdIndex; wire[4:0] rs1Index; wire[4:0] rs2Index;
	wire[2:0] funct3; wire[6:0] funct7;
	wire isCompressed;
	wire isLUI; wire isAUIPC; wire isJAL; wire isJALR; wire isBranch; wire isLoad; wire isStore;
	wire isALUImmBase; wire isALUImmNormal; wire isALUImmShift; wire isALUImm; wire isALU;
	wire isSystem; 
	wire isCSR; wire isCSRIMM; wire isCSRRW; wire isCSRRS; wire isCSRRC; 
	InstructionDecode decode(
		.currentInstruction(currentInstruction),
		.isNOP(pipeStall),
		.opcode(opcode),
		.rdIndex(rdIndex), .rs1Index(rs1Index), .rs2Index(rs2Index),
		.funct3(funct3), .funct7(funct7),
		.isCompressed(isCompressed),
		.isLUI(isLUI), .isAUIPC(isAUIPC), .isJAL(isJAL), .isJALR(isJALR), .isBranch(isBranch), .isLoad(isLoad), .isStore(isStore),
		.isALUImmBase(isALUImmBase), .isALUImmNormal(isALUImmNormal), .isALUImmShift(isALUImmShift), .isALUImm(isALUImm), .isALU(isALU),
		.isFence(isFence), .isSystem(isSystem),
		.isCSR(isCSR), .isCSRIMM(isCSRIMM), .isCSRRW(isCSRRW), .isCSRRS(isCSRRS), .isCSRRC(isCSRRC),
		.isECALL(isECALL), .isEBREAK(isEBREAK), .isRET(isRET),
		.invalidInstruction(invalidInstruction)
	);

	// Immediate Decode
	wire[31:0] imm_I = {currentInstruction[31] ? 21'h1F_FFFF : 21'h00_0000, currentInstruction[30:25], currentInstruction[24:21], currentInstruction[20]};
	wire[31:0] imm_S = {currentInstruction[31] ? 21'h1F_FFFF : 21'h00_0000, currentInstruction[30:25], currentInstruction[11:8] , currentInstruction[7]};
	wire[31:0] imm_B = {currentInstruction[31] ? 20'hF_FFFF  : 20'h0_0000 , currentInstruction[7]    , currentInstruction[30:25], currentInstruction[11:8] , 1'b0};
	wire[31:0] imm_U = {currentInstruction[31]							  , currentInstruction[30:20], currentInstruction[19:12], 12'h000};
	wire[31:0] imm_J = {currentInstruction[31] ? 12'hFFF : 12'h000 		  , currentInstruction[19:12], currentInstruction[20]	, currentInstruction[30:25], currentInstruction[24:21], 1'b0};


	// Setup inputs for ALU and branch control
	wire[31:0] inputA = isAUIPC ? programCounter : rs1Data;
	reg[31:0] inputB;
	always @(*) begin
		case (1'b1)
			isAUIPC : inputB <= imm_U;
			isALUImm: inputB <= imm_I;
			isLoad 	: inputB <= imm_I;
			isStore : inputB <= imm_S;
			default: inputB <= rs2Data;
		endcase
	end

	// The use of A-B for comparison is based on https://github.com/BrunoLevy/learn-fpga/tree/master/FemtoRV/TUTORIALS/FROM_BLINKER_TO_RISCV#from-blinker-to-risc-v
	wire[31:0] aluAPlusB = inputA + inputB;
	wire[32:0] aluACompareB = { 1'b0, inputA } - { 1'b0, inputB };
	wire[31:0] aluAMinusB = aluACompareB[31:0];
	wire aluAEqualsB = aluAMinusB == 32'b0;
	wire aluALessThanB = inputA[31] ^ inputB[31] ? inputA[31] : aluACompareB[32];
	wire aluALessThanBUnsigned = aluACompareB[32];

	// Jump and branch control
	reg takeBranch;
	always @(*) begin
		if (isBranch) begin
			case (funct3)
				/*BEQ*/  3'b000: takeBranch <= aluAEqualsB;
				/*BNE*/  3'b001: takeBranch <= !aluAEqualsB;
				//*None*/ 3'b010: takeBranch <= 1'b0;
				//*None*/ 3'b011: takeBranch <= 1'b0;
				/*BLT*/  3'b100: takeBranch <= aluALessThanB;
				/*BGE*/  3'b101: takeBranch <= !aluALessThanB;
				/*BLTU*/ 3'b110: takeBranch <= aluALessThanBUnsigned;
				/*BGEU*/ 3'b111: takeBranch <= !aluALessThanBUnsigned;
						default: takeBranch <= 1'b0;
			endcase
		end else begin
			takeBranch <= 1'b0;
		end
	end

	wire[31:0] programCounterLink = programCounter + (isCompressed ? 2 : 4);

	reg[31:0] nextProgramCounterBase;
	always @(*) begin
		case (1'b1)
			isJAL 	   : nextProgramCounterBase <= programCounter;
			isJALR     : nextProgramCounterBase <= rs1Data;
			takeBranch : nextProgramCounterBase <= programCounter;
			default    : nextProgramCounterBase <= programCounterLink;
		endcase
	end

	reg[31:0] nextProgramCounterOffset;
	always @(*) begin
		case (1'b1)
			isJAL 	   : nextProgramCounterOffset <= imm_J;
			isJALR     : nextProgramCounterOffset <= imm_I;
			takeBranch : nextProgramCounterOffset <= imm_B;
			default    : nextProgramCounterOffset <= 32'b0;
		endcase
	end

	wire[31:0] nextProgramCounterWord = nextProgramCounterBase + nextProgramCounterOffset;
	wire[31:0] nextProgramCounterCompressed = programCounterLink; // TODO: Need to implement compressed branch and jump instructions
	wire[31:0] nextProgramCounterFull = isCompressed ? nextProgramCounterCompressed : nextProgramCounterWord;
	assign isJump = isJAL || isJALR || isBranch;
	assign jumpEnable = isJAL || isJALR || takeBranch;
	assign failedBranch = isBranch && !takeBranch;
	assign nextProgramCounter = { nextProgramCounterFull[31:1] , 1'b0};
	assign jumpMissaligned = !isCompressed && |nextProgramCounter[1:0] && (isJAL || isJALR || takeBranch);

	// ALU	
	wire aluAlt = funct7 == 7'b0100000 && (isALU || isALUImmShift);
	
	// Using only a single shifter also from https://github.com/BrunoLevy/learn-fpga/tree/master/FemtoRV/TUTORIALS/FROM_BLINKER_TO_RISCV#from-blinker-to-risc-v
	// Although I feel like there is an easier way to flip bit orderings
	function [31:0] flipBits32 (input [31:0] x);
		flipBits32 = { x[ 0], x[ 1], x[ 2], x[ 3], x[ 4], x[ 5], x[ 6], x[ 7], 
					   x[ 8], x[ 9], x[10], x[11], x[12], x[13], x[14], x[15], 
					   x[16], x[17], x[18], x[19], x[20], x[21], x[22], x[23],
					   x[24], x[25], x[26], x[27], x[28], x[29], x[30], x[31] };
	endfunction

	wire isLeftShift = funct3 == 3'b001;
	wire[31:0] shiftInput = isLeftShift ? flipBits32(inputA) : inputA;
	wire signed[32:0] signedShiftInput = { aluAlt && shiftInput[31] && !isLeftShift, shiftInput };
	wire[32:0] aluShifter = $signed(signedShiftInput >>> inputB[4:0]);
	wire[31:0] rightShift = aluShifter[31:0];
	wire[31:0] leftShift = flipBits32(rightShift);

	reg[31:0] aluValue;
	always @(*) begin
		case (funct3)
			/*ADD*/  3'b000: aluValue <= aluAlt ? aluAMinusB : aluAPlusB;
			/*SLL*/  3'b001: aluValue <= leftShift;
			/*SLT*/  3'b010: aluValue <= {31'b0, aluALessThanB};
			/*SLTU*/ 3'b011: aluValue <= {31'b0, aluALessThanBUnsigned};
			/*XOR*/  3'b100: aluValue <= inputA ^ inputB;
			/*SRL*/  3'b101: aluValue <= rightShift;
			/*OR*/   3'b110: aluValue <= inputA | inputB;
			/*AND*/  3'b111: aluValue <= inputA & inputB;
					default: aluValue <= 32'b0;
		endcase
	end

	wire[31:0] csrRS1Data = isCSRIMM ? { 27'b0, rs1Index} : rs1Data;

	reg[31:0] csrWriteData;
	always @(*) begin
		if (isCSR) begin			
			if (isCSRRW) csrWriteData <= csrRS1Data;
			else if (isCSRRS) csrWriteData <= csrReadData | csrRS1Data;
			else if (isCSRRC) csrWriteData <= csrReadData & ~csrRS1Data;
			else csrWriteData <= 32'b0;
		end else begin
			csrWriteData <= 32'b0;
		end 
	end

	wire csrRead = isCSRRC || isCSRRS || (isCSR && |rdIndex);
	wire needStore = isLUI || isAUIPC || isJAL || isJALR || isALU || isALUImm || isLoad || csrRead;

	reg[31:0] currentData;
	always @(*) begin
		case (1'b1)
			isLUI			   : currentData <= imm_U;
			isAUIPC			   : currentData <= aluAPlusB;
			isJAL			   : currentData <= programCounterLink;
			isJALR	   		   : currentData <= programCounterLink;
			(isALU || isALUImm): currentData <= aluValue;
			isLoad 			   : currentData <= aluAPlusB;
			csrRead	   		   : currentData <= csrWriteData;
			default: currentData <= 32'b0;
		endcase
	end

	// Memory interface
	wire[31:0] targetMemoryAddress = aluAPlusB;
	wire loadSigned    = (funct3 == 3'b000) || (funct3 == 3'b001);
	wire loadStoreByte = funct3[1:0] == 2'b00;
	wire loadStoreHalf = funct3[1:0] == 2'b01;
	wire loadStoreWord = funct3 == 3'b010;
	reg[3:0] baseByteMask;
	always @(*) begin
		if ((isLoad || isStore)) begin
			if (loadStoreWord) baseByteMask <= 4'b1111;
			else if (loadStoreHalf) baseByteMask <= 4'b0011;
			else if (loadStoreByte) baseByteMask <= 4'b0001;
			else baseByteMask <= 4'b0000;
		end else begin
			baseByteMask <= 4'b0000;
		end
	end

	wire[6:0] loadStoreByteMask = {3'b0, baseByteMask} << targetMemoryAddress[1:0];
	wire loadStoreByteMaskValid = |(loadStoreByteMask[3:0]);
	wire isAddressMisaligned = |loadStoreByteMask[6:4] || (loadStoreHalf && targetMemoryAddress[1:0] == 2'h1);
	assign fullMemoryAddress = targetMemoryAddress;
	assign addressMisaligned_load = isAddressMisaligned && isLoad;
	assign addressMisaligned_store = isAddressMisaligned && isStore;
	wire shouldLoad  = loadStoreByteMaskValid && !isAddressMisaligned && isLoad;
	wire shouldStore = loadStoreByteMaskValid && !isAddressMisaligned && isStore;
	wire shouldLoadOrStore = shouldLoad || shouldStore;

	reg[31:0] dataOut;
	always @(*) begin
		case (targetMemoryAddress[1:0])
			2'b00: dataOut = {
					baseByteMask[3] ? rs2Data[31:24] : 8'h00,
					baseByteMask[2] ? rs2Data[23:16] : 8'h00,
					baseByteMask[1] ? rs2Data[15:8]  : 8'h00,
					baseByteMask[0] ? rs2Data[7:0]   : 8'h00
				};

			2'b01: dataOut = {
					baseByteMask[2] ? rs2Data[23:16] : 8'h00,
					baseByteMask[1] ? rs2Data[15:8]  : 8'h00,
					baseByteMask[0] ? rs2Data[7:0]   : 8'h00,
					8'h00
				};

			2'b10: dataOut = {
					baseByteMask[1] ? rs2Data[15:8]  : 8'h00,
					baseByteMask[0] ? rs2Data[7:0]   : 8'h00,
					8'h00,
					8'h00
				};

			2'b11: dataOut = {
					baseByteMask[0] ? rs2Data[7:0]   : 8'h00,
					8'h00,
					8'h00,
					8'h00
				};
		endcase
	end

	// Register read control
	assign rs1Address = rs1Index;
	assign rs2Address = rs2Index;

	// CSR read control
	assign csrReadAddress = currentInstruction[31:20];
	assign csrReadEnable = csrRead && !pipeStall;

	// Result register control
	assign operationResultStoreEnable = needStore && !pipeStall;
	assign operationResult = currentData;

	// Load/Store control
	assign memoryEnable = shouldLoadOrStore && !pipeStall;
	assign memoryWriteEnable = shouldStore && !pipeStall;
	assign memoryByteSelect = shouldLoadOrStore ? loadStoreByteMask[3:0] : 4'b0000;
	assign memoryAddress = shouldLoadOrStore ? { targetMemoryAddress[31:2], 2'b00 } : 32'b0;
	assign memoryWriteData = dataOut;

endmodulemodule PipeStage (
		input wire clk,
		input wire rst,

		// Pipe control
		input wire stepPipe,
		input wire pipeStall,
		output reg currentPipeStall,
		output wire active,
		input wire[31:0] currentInstruction,
		output reg[31:0] lastInstruction
	);

	always @(posedge clk) begin
		if (rst) begin
			currentPipeStall <= 1'b1;
			lastInstruction <= 32'b0;
		end else begin
			if (stepPipe) begin
				currentPipeStall <= pipeStall;
				if (!pipeStall) lastInstruction <= currentInstruction;
			end
		end
	end

	assign active = !pipeStall;
	
endmodulemodule PipeStore (
		input wire clk,
		input wire rst,

		// Pipe control
		input wire stepPipe,
		input wire pipeStall,
		output wire currentPipeStall,
		output wire active,
		input wire[31:0] currentInstruction,
		output wire[31:0] lastInstruction,
		output wire invalidInstruction,

		// Memory control
		output wire expectingLoad,

		// Store inputs
		input wire[31:0] memoryDataRead,
		input wire[31:0] aluResultData,
		input wire[31:0] csrData,

		// Register store control
		output wire[4:0] registerWriteAddress,
		output wire[31:0] registerWriteData,
		output wire registerWriteEnable,

		// CSR store control
		output wire[11:0] csrWriteAddress,
		output wire[31:0] csrWriteData,
		output wire csrWriteEnable,

		// Stall control
		output wire isJump,
		output wire isFence,
		output wire isRET
	);
	
	// Pipe control
	PipeStage pipeStage(
		.clk(clk),
		.rst(rst),
		.stepPipe(stepPipe),
		.pipeStall(pipeStall),
		.currentPipeStall(currentPipeStall),
		.active(active),
		.currentInstruction(currentInstruction),
		.lastInstruction(lastInstruction));

	// Instruction decode
	wire[6:0] opcode;
	wire[4:0] rdIndex; wire[4:0] rs1Index; wire[4:0] rs2Index;
	wire[2:0] funct3; wire[6:0] funct7;
	wire isCompressed;
	wire isLUI; wire isAUIPC; wire isJAL; wire isJALR; wire isBranch; wire isLoad; wire isStore;
	wire isALUImmBase; wire isALUImmNormal; wire isALUImmShift; wire isALUImm; wire isALU;
	wire isSystem; 
	wire isCSR; wire isCSRIMM; wire isCSRRW; wire isCSRRS; wire isCSRRC; 
	wire isECALL; wire isEBREAK;
	InstructionDecode decode(
		.currentInstruction(currentInstruction),
		.isNOP(pipeStall),
		.opcode(opcode),
		.rdIndex(rdIndex), .rs1Index(rs1Index), .rs2Index(rs2Index),
		.funct3(funct3), .funct7(funct7),
		.isCompressed(isCompressed),
		.isLUI(isLUI), .isAUIPC(isAUIPC), .isJAL(isJAL), .isJALR(isJALR), .isBranch(isBranch), .isLoad(isLoad), .isStore(isStore),
		.isALUImmBase(isALUImmBase), .isALUImmNormal(isALUImmNormal), .isALUImmShift(isALUImmShift), .isALUImm(isALUImm), .isALU(isALU),
		.isFence(isFence), .isSystem(isSystem),
		.isCSR(isCSR), .isCSRIMM(isCSRIMM), .isCSRRW(isCSRRW), .isCSRRS(isCSRRS), .isCSRRC(isCSRRC),
		.isECALL(isECALL), .isEBREAK(isEBREAK), .isRET(isRET),
		.invalidInstruction(invalidInstruction)
	);

	// Memory connections
	wire[31:0] targetMemoryAddress = aluResultData;
	wire loadSigned    = (funct3 == 3'b000) || (funct3 == 3'b001);
	wire loadStoreByte = funct3[1:0] == 2'b00;
	wire loadStoreHalf = funct3[1:0] == 2'b01;
	wire loadStoreWord = funct3 == 3'b010;
	reg[3:0] baseByteMask;
	always @(*) begin
		if (isLoad || isStore) begin
			if (loadStoreWord) baseByteMask <= 4'b1111;
			else if (loadStoreHalf) baseByteMask <= 4'b0011;
			else if (loadStoreByte) baseByteMask <= 4'b0001;
			else baseByteMask <= 4'b0000;
		end else begin
			baseByteMask <= 4'b0000;
		end
	end

	reg signExtend;
	always @(*) begin
		if (loadSigned) begin
			if (loadStoreByte) begin
				case (targetMemoryAddress[1:0])
					2'b00: signExtend <= memoryDataRead[7];
					2'b01: signExtend <= memoryDataRead[15];
					2'b10: signExtend <= memoryDataRead[23];
					2'b11: signExtend <= memoryDataRead[31];
				endcase
			end else if (loadStoreHalf) begin
				case (targetMemoryAddress[1:0])
					2'b00: signExtend <= memoryDataRead[15];
					2'b01: signExtend <= memoryDataRead[23];
					2'b10: signExtend <= memoryDataRead[31];
					2'b11: signExtend <= 1'b0;
				endcase
			end else begin
				signExtend <= 1'b0;
			end
		end else begin
			signExtend <= 1'b0;
		end
	end

	wire[7:0] signExtendByte = signExtend ? 8'hFF : 8'h00;

	wire[6:0] loadStoreByteMask = {3'b0, baseByteMask} << targetMemoryAddress[1:0];
	wire loadStoreByteMaskValid = |(loadStoreByteMask[3:0]);
	wire addressMissaligned = |loadStoreByteMask[6:4];
	wire shouldLoad  = loadStoreByteMaskValid && !addressMissaligned && isLoad;

	reg[31:0] dataIn;
	always @(*) begin
		case (targetMemoryAddress[1:0])
			2'b00: dataIn = {
					loadStoreByteMask[3] ? memoryDataRead[31:24] : signExtendByte,
					loadStoreByteMask[2] ? memoryDataRead[23:16] : signExtendByte,
					loadStoreByteMask[1] ? memoryDataRead[15:8]  : signExtendByte,
					loadStoreByteMask[0] ? memoryDataRead[7:0]   : 8'h00
				};

			2'b01: dataIn = {
					signExtendByte,
					loadStoreByteMask[3] ? memoryDataRead[31:24] : signExtendByte,
					loadStoreByteMask[2] ? memoryDataRead[23:16] : signExtendByte,
					loadStoreByteMask[1] ? memoryDataRead[15:8]  : 8'h00
				};

			2'b10: dataIn = {
					signExtendByte,
					signExtendByte,
					loadStoreByteMask[3] ? memoryDataRead[31:24] : signExtendByte,
					loadStoreByteMask[2] ? memoryDataRead[23:16] : 8'h00
				};

			2'b11: dataIn = {
					signExtendByte,
					signExtendByte,
					signExtendByte,
					loadStoreByteMask[3] ? memoryDataRead[31:24] : 8'h00
				};
		endcase
	end

	// Register Write
	wire csrWrite = isCSRRW || (isCSR && |rdIndex);
	wire integerRegisterWriteEn = isLUI || isAUIPC || isJAL || isJALR || isALU || isALUImm || isLoad || csrWrite;
	reg[31:0] integerRegisterWriteData;
	always @(*) begin
		case (1'b1)
			isLUI			   : integerRegisterWriteData <= aluResultData;
			isAUIPC			   : integerRegisterWriteData <= aluResultData;
			isJAL			   : integerRegisterWriteData <= aluResultData;
			isJALR	   		   : integerRegisterWriteData <= aluResultData;
			shouldLoad  	   : integerRegisterWriteData <= dataIn;
			(isALU || isALUImm): integerRegisterWriteData <= aluResultData;
			csrWrite   		   : integerRegisterWriteData <= csrData;
			default: integerRegisterWriteData <= 32'b0;
		endcase
	end

	// Memory control
	assign expectingLoad = shouldLoad;
	
	// Register write control
	assign registerWriteAddress = rdIndex;
	assign registerWriteData = integerRegisterWriteData;
	assign registerWriteEnable = integerRegisterWriteEn && !pipeStall;

	// CSR write control
	assign csrWriteAddress = currentInstruction[31:20];
	assign csrWriteData = aluResultData;
	assign csrWriteEnable = csrWrite && !pipeStall;

	// Stall control
	assign isJump = isJAL || isJALR || isBranch;

endmodulemodule InstructionDecode (
		input wire[31:0] currentInstruction,
		input wire isNOP,
		output reg[6:0] opcode,
		output reg[4:0] rdIndex,
		output reg[4:0] rs1Index,
		output reg[4:0] rs2Index,
		output reg[2:0] funct3,
		output reg[6:0] funct7,
		output reg isCompressed,
		output reg isLUI,
		output reg isAUIPC,
		output reg isJAL,
		output reg isJALR,
		output reg isBranch,
		output reg isLoad,
		output reg isStore,
		output reg isALUImmBase,
		output reg isALUImmNormal,
		output reg isALUImmShift,
		output reg isALUImm,
		output reg isALU,
		output reg isFence,
		output reg isSystem,
		output reg isCSR,
		output reg isCSRIMM,
		output reg isCSRRW,
		output reg isCSRRS,
		output reg isCSRRC,
		output reg isECALL,
		output reg isEBREAK,
		output reg isRET,
		output reg invalidInstruction
	);
	
	

	// Instruction decode
	always @(*) begin
		if (isNOP) begin
			opcode <= 7'b0;
			rdIndex <= 5'b0;
			rs1Index <= 5'b0;
			rs2Index <= 5'b0;
			funct3 <= 3'b0;
			funct7 <= 7'b0;
			isCompressed <= 1'b0;
		end else begin
			opcode <= currentInstruction[6:0];
			rdIndex <= currentInstruction[11:7];
			rs1Index <= currentInstruction[19:15];
			rs2Index <= currentInstruction[24:20];
			funct3 <= currentInstruction[14:12];
			funct7 <= currentInstruction[31:25];
			isCompressed <= opcode[1:0] != 2'b11;
		end
	end

	// Instruction decode
	always @(*) begin
		if (isNOP) begin
			isLUI 		   <= 1'b0;
			isAUIPC 	   <= 1'b0;
			isJAL 		   <= 1'b0;
			isJALR   	   <= 1'b0;
			isBranch 	   <= 1'b0;
			isLoad   	   <= 1'b0;
			isStore  	   <= 1'b0;
			isALUImmBase   <= 1'b0;
			isALUImmNormal <= 1'b0;
			isALUImmShift  <= 1'b0;
			isALUImm 	   <= 1'b0;
			isALU 	 	   <= 1'b0;
			isFence  	   <= 1'b0;
			isSystem 	   <= 1'b0;
		end else begin
			isLUI 		   <= (opcode == 7'b0110111);
			isAUIPC 	   <= (opcode == 7'b0010111);
			isJAL 		   <= (opcode == 7'b1101111);
			isJALR   	   <= (opcode == 7'b1100111) && (funct3 == 3'b000);
			isBranch 	   <= (opcode == 7'b1100011) && (funct3 != 3'b010) && (funct3 != 3'b011);
			isLoad   	   <= (opcode == 7'b0000011) && (funct3 == 3'b000 || funct3 == 3'b001 || funct3 == 3'b010 || funct3 == 3'b100 || funct3 == 3'b101);
			isStore  	   <= (opcode == 7'b0100011) && (funct3 == 3'b000 || funct3 == 3'b001 || funct3 == 3'b010);
			isALUImmBase   <= (opcode == 7'b0010011);
			isALUImmNormal <= isALUImmBase && funct3 != 3'b001 && funct3 != 3'b101;
			isALUImmShift  <= isALUImmBase && ((funct3 == 3'b001 && funct7 == 7'b0000000) || (funct3 == 3'b101 && (funct7 == 7'b0000000 || funct7 == 7'b0100000)));
			isALUImm 	   <= isALUImmShift || isALUImmNormal;
			isALU 	 	   <= (opcode == 7'b0110011) && (funct7 == 7'b0000000 || ((funct7 == 7'b0100000) && (funct3 == 3'b000 || funct3 == 3'b101)));
			isFence  	   <= (opcode == 7'b0001111) && (funct3 == 3'b000);
			isSystem 	   <= (opcode == 7'b1110011);
		end
	end
	
	
	// System commands
	always @(*) begin
		if (isNOP) begin
			isCSR 	 <= 1'b0;
			isCSRIMM <= 1'b0;
			isCSRRW  <= 1'b0;
			isCSRRS  <= 1'b0;
			isCSRRC  <= 1'b0;
			isECALL  <= 1'b0;
			isEBREAK <= 1'b0;
			isRET 	 <= 1'b0;
		end else begin
			isCSR 	 <= isSystem && (funct3 != 3'b000);
			isCSRIMM <= isCSR && funct3[2];
			isCSRRW  <= isCSR && (funct3[1:0] == 2'b01);
			isCSRRS  <= isCSR && (funct3[1:0] == 2'b10);
			isCSRRC  <= isCSR && (funct3[1:0] == 2'b11);
			isECALL  <= isSystem && (currentInstruction[31:7] == 25'b0000000000000000000000000);
			isEBREAK <= isSystem && (currentInstruction[31:7] == 25'b0000000000010000000000000);
			isRET 	 <= isSystem && (currentInstruction[31:7] == 25'b0011000000100000000000000);
		end
	end

	wire validSystemCommand = isCSR || isECALL || isEBREAK || isRET;

	always @(*) begin
		if (isNOP) begin
			invalidInstruction <= 1'b0;
		end else begin
			case ({ isLUI, isAUIPC, isJAL, isJALR, isBranch, isLoad, isStore, isALUImm, isALU, isFence, isSystem })
				'b00000000001: invalidInstruction <= 1'b0;
				'b00000000010: invalidInstruction <= 1'b0;
				'b00000000100: invalidInstruction <= 1'b0;
				'b00000001000: invalidInstruction <= 1'b0;
				'b00000010000: invalidInstruction <= 1'b0;
				'b00000100000: invalidInstruction <= 1'b0;
				'b00001000000: invalidInstruction <= 1'b0;
				'b00010000000: invalidInstruction <= 1'b0;
				'b00100000000: invalidInstruction <= 1'b0;
				'b01000000000: invalidInstruction <= 1'b0;
				'b10000000000: invalidInstruction <= validSystemCommand;
				default: invalidInstruction <= 1'b1;
			endcase
		end
	end

endmodulemodule MisalignedMemoryController (
		input wire clk,
		input wire rst,

		// External memory interface
		output wire[31:0] external_memoryAddress,
		output wire[3:0] external_memoryByteSelect,
		output wire external_memoryWriteEnable,
		output wire external_memoryReadEnable,
		output wire[31:0] external_memoryDataWrite,
		input wire[31:0] external_memoryDataRead,
		input wire external_memoryBusy,
		input wire external_memoryAccessFault,
		input wire external_addressBreakpoint,
		
		// Internal memory interface
		output wire[31:0] internal_memoryAddress,
		output wire[3:0] internal_memoryByteSelect,
		output wire internal_memoryWriteEnable,
		output wire internal_memoryReadEnable,
		output wire[31:0] internal_memoryDataWrite,
		input wire[31:0] internal_memoryDataRead,
		input wire internal_memoryBusy,
		input wire internal_memoryAccessFault,
		input wire internal_addressBreakpoint
	);
	


endmodulemodule CSR (
		input wire clk,
		input wire rst,

		// CSR interface
		input wire csrWriteEnable,
		input wire csrReadEnable,
		input wire[11:0] csrWriteAddress,
		input wire[11:0] csrReadAddress,
		input wire[31:0] csrWriteData,
		output reg[31:0] csrReadData,

		// System interface
		input wire[7:0] coreIndex,
		input wire[10:0] manufacturerID,
		input wire[15:0] partID,
		input wire[3:0] versionID,
		input wire[25:0] extensions,
		input wire instructionCompleted,

		// System trap interface
		input wire[31:0] programCounter,
		input wire[31:0] currentInstruction,
		input wire[31:0] instruction_memoryAddress,
		input wire[31:0] data_memoryAddress,
		input wire isMachineTimerInterrupt,
		input wire isMachineExternalInterrupt,
		input wire isMachineSoftwareInterrupt,
		input wire isFetchAddressMisaligned,
		input wire isDataAddressMisaligned_load,
		input wire isDataAddressMisaligned_store,
		input wire isJumpMissaligned,
		input wire isFetchAccessFault,
		input wire isDataAccessFault_load,
		input wire isDataAccessFault_store,
		input wire isInvalidInstruction,
		input wire isEBREAK,
		input wire isECALL,
		input wire isFetchAddressBreakpoint,
		input wire isDataAddressBreakpoint,
		input wire[15:0] userInterrupts,
		input wire trapReturn,
		output wire inTrap,
		output wire[31:0] trapVector,
		output wire[31:0] trapReturnVector
	);

	// Cylce
	wire[63:0] cycleCount;
	wire[31:0] cycleTimerReadData;
	wire cycleTimerRequestOutput;
	CSR_TimerRegister #(.ADDRESS_LOWER(12'hC00), .ADDRESS_UPPER(12'hC80)) cycleTimer (
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(cycleTimerReadData),
		.csrRequestOutput(cycleTimerRequestOutput),
		.count(1'b1),
		.value(cycleCount));

	// Time
	// Time register is duplicate of cycle register
	wire[31:0] timeTimerReadDataLower;
	wire timeTimerRequestOutputLower;
	CSR_ReadRegister #(.ADDRESS(12'hC01)) timeTimerLower(
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(timeTimerReadDataLower),
		.csrRequestOutput(timeTimerRequestOutputLower),
		.value(cycleCount[31:0]));

	wire[31:0] timeTimerReadDataUpper;
	wire timeTimerRequestOutputUpper;
	CSR_ReadRegister #(.ADDRESS(12'hC81)) timeTimerUpper(
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(timeTimerReadDataUpper),
		.csrRequestOutput(timeTimerRequestOutputUpper),
		.value(cycleCount[63:32]));

	// Instret
	wire[31:0] instretTimerReadData;
	wire instretTimerRequestOutput;
	CSR_TimerRegister #(.ADDRESS_LOWER(12'hC02), .ADDRESS_UPPER(12'hC82)) instretTimer (
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(instretTimerReadData),
		.csrRequestOutput(instretTimerRequestOutput),
		.count(instructionCompleted));

	// Vendor ID
	wire[31:0] vendorIDReadData;
	wire vendorIDRequestOutput;
	CSR_ReadRegister #(.ADDRESS(12'hF11)) vendorID(
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(vendorIDReadData),
		.csrRequestOutput(vendorIDRequestOutput),
		.value({ 21'b0, manufacturerID }));

	// Architecture ID
	wire[31:0] archIDReadData;
	wire archIDRequestOutput;
	CSR_ReadRegister #(.ADDRESS(12'hF12)) archID(
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(archIDReadData),
		.csrRequestOutput(archIDRequestOutput),
		.value({ 16'b0, partID }));

	// Implementation ID
	wire[31:0] implIDReadData;
	wire implIDRequestOutput;
	CSR_ReadRegister #(.ADDRESS(12'hF13)) implID(
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(implIDReadData),
		.csrRequestOutput(implIDRequestOutput),
		.value({ 28'b0, versionID }));

	// Hardware thread ID
	wire[31:0] coreIDReadData;
	wire coreIDRequestOutput;
	CSR_ReadRegister #(.ADDRESS(12'hF14)) coreID(
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(coreIDReadData),
		.csrRequestOutput(coreIDRequestOutput),
		.value({ 24'b0, coreIndex }));

	// Pointer to configuration data structure
	wire[31:0] configPointerReadData;
	wire configPointerRequestOutput;
	wire[31:0] configPointerValue_nc;
	CSR_ConfigurationRegister #(.ADDRESS(12'hF15)) mconfigptr(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(configPointerReadData),
		.csrRequestOutput(configPointerRequestOutput),
		.value(configPointerValue_nc));

	// ISA
	wire[31:0] misaReadData;
	wire misaRequestOutput;
	CSR_ReadRegister #(.ADDRESS(12'h301)) misa(
		.clk(clk),
		.rst(rst),
		.csrReadEnable(csrReadEnable),
		.csrReadAddress(csrReadAddress),
		.csrReadData(misaReadData),
		.csrRequestOutput(misaRequestOutput),
		.value({ 2'b01, 4'b0, extensions }));

	// Trap handling
	wire[31:0] trapsReadData;
	wire trapsRequestOutput;
	Traps traps(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(trapsReadData),
		.requestOutput(trapsRequestOutput),
		.programCounter(programCounter),
		.currentInstruction(currentInstruction),
		.instruction_memoryAddress(instruction_memoryAddress),
		.data_memoryAddress(data_memoryAddress),
		.isMachineTimerInterrupt(isMachineTimerInterrupt),
		.isMachineExternalInterrupt(isMachineExternalInterrupt),
		.isMachineSoftwareInterrupt(isMachineSoftwareInterrupt),
		.isFetchAddressMisaligned(isFetchAddressMisaligned),
		.isDataAddressMisaligned_load(isDataAddressMisaligned_load),
		.isDataAddressMisaligned_store(isDataAddressMisaligned_store),
		.isJumpMissaligned(isJumpMissaligned),
		.isFetchAccessFault(isFetchAccessFault),
		.isDataAccessFault_load(isDataAccessFault_load),
		.isDataAccessFault_store(isDataAccessFault_store),
		.isInvalidInstruction(isInvalidInstruction),
		.isEBREAK(isEBREAK),
		.isECALL(isECALL),
		.isFetchAddressBreakpoint(isFetchAddressBreakpoint),
		.isDataAddressBreakpoint(isDataAddressBreakpoint),
		.userInterrupts(userInterrupts),
		.trapReturn(trapReturn),
		.inTrap(inTrap),
		.trapVector(trapVector),
		.trapReturnVector(trapReturnVector));

	always @(*) begin
		case (1'b1)
			// Timers
			cycleTimerRequestOutput: csrReadData <= cycleTimerReadData;
			timeTimerRequestOutputLower: csrReadData <= timeTimerReadDataLower;
			timeTimerRequestOutputUpper: csrReadData <= timeTimerReadDataUpper;
			instretTimerRequestOutput: csrReadData <= instretTimerReadData;
			
			// Machine info
			vendorIDRequestOutput: csrReadData <= vendorIDReadData;
			archIDRequestOutput: csrReadData <= archIDReadData;
			implIDRequestOutput: csrReadData <= implIDReadData;
			coreIDRequestOutput: csrReadData <= coreIDReadData;
			configPointerRequestOutput: csrReadData <= configPointerReadData;
			misaRequestOutput: csrReadData <= misaReadData;

			// Traps
			trapsRequestOutput: csrReadData <= trapsReadData;

			default: csrReadData <= 32'b0;
		endcase
	end

endmodulemodule CSR_ConfigurationRegister #(
		parameter ADDRESS = 12'h000,
		parameter DEFAULT = 32'b0
	)(
		input wire clk,
		input wire rst,

		// CSR interface
		input wire csrWriteEnable,
		input wire csrReadEnable,
		input wire[11:0] csrWriteAddress,
		input wire[11:0] csrReadAddress,
		input wire[31:0] csrWriteData,
		output wire[31:0] csrReadData,
		output wire csrRequestOutput,

		// System interface
		output wire[31:0] value
	);
	
	wire csrWriteEnabled = csrWriteAddress == ADDRESS;
	wire csrReadEnabled = csrReadAddress == ADDRESS;

	reg[31:0] currentValue = DEFAULT;

	always @(posedge clk) begin
		if (rst) begin
			currentValue <= DEFAULT;
		end else begin
			if (csrWriteEnabled && csrWriteEnable) currentValue <= csrWriteData;
		end
	end

	assign csrReadData = csrReadEnabled && csrReadEnable ? currentValue : 32'b0;
	assign csrRequestOutput = csrReadEnabled && csrReadEnable;

	assign value = currentValue;
	
endmodulemodule CSR_DataRegister #(
		parameter ADDRESS = 12'h000
	)(
		input wire clk,
		input wire rst,

		// CSR interface
		input wire csrWriteEnable,
		input wire csrReadEnable,
		input wire[11:0] csrWriteAddress,
		input wire[11:0] csrReadAddress,
		input wire[31:0] csrWriteData,
		output wire[31:0] csrReadData,
		output wire csrRequestOutput,

		// System interface
		input wire[31:0] readData,
		output wire readDataEnable,
		output wire[31:0] writeData,
		output wire writeDataEnable
	);
	
	wire csrWriteEnabled = csrWriteAddress == ADDRESS;
	wire csrReadEnabled = csrReadAddress == ADDRESS;

	assign csrReadData = csrReadEnabled && csrReadEnable ? readData : 32'b0;
	assign readDataEnable = csrReadEnabled && csrReadEnable;
	assign writeData = csrWriteData;
	assign writeDataEnable = csrWriteEnabled && csrWriteEnable;

	assign csrRequestOutput = csrReadEnabled && csrReadEnable;
	
endmodulemodule CSR_ReadRegister #(
		parameter ADDRESS = 12'h000
	)(
		input wire clk,
		input wire rst,

		// CSR interface
		input wire csrReadEnable,
		input wire[11:0] csrReadAddress,
		output wire[31:0] csrReadData,
		output wire csrRequestOutput,

		// System interface
		input wire[31:0] value
	);
	
	wire csrReadEnabled = csrReadAddress == ADDRESS;

	assign csrReadData = csrReadEnabled && csrReadEnable ? value : 32'b0;
	assign csrRequestOutput = csrReadEnabled && csrReadEnable;

endmodulemodule CSR_TimerRegister #(
		parameter ADDRESS_LOWER = 12'h000,
		parameter ADDRESS_UPPER = 12'h000
	)(
		input wire clk,
		input wire rst,

		// CSR interface
		input wire csrReadEnable,
		input wire[11:0] csrReadAddress,
		output reg[31:0] csrReadData,
		output wire csrRequestOutput,

		// System interface
		input wire count,
		output wire[63:0] value
	);
	
	wire csrReadEnabledLower = csrReadAddress == ADDRESS_LOWER;
	wire csrReadEnabledUpper = csrReadAddress == ADDRESS_UPPER;

	reg[63:0] currentValue = 64'b0;

	always @(posedge clk) begin
		if (rst) begin
			currentValue <= 64'b0;
		end else begin
			if (count) currentValue <= currentValue + 1;
		end
	end

	always @(*) begin
		if (csrReadEnable) begin
			if (csrReadEnabledLower) csrReadData <= currentValue[31:0];
			else if (csrReadEnabledUpper) csrReadData <= currentValue[63:32];
			else csrReadData <= 32'b0;
		end else begin
			csrReadData <= 32'b0;
		end 
	end

	assign csrRequestOutput = (csrReadEnabledLower || csrReadEnabledUpper) && csrReadEnable;
	
	assign value = currentValue;
	
endmodulemodule Traps (
		input wire clk,
		input wire rst,

		// CSR interface
		input wire csrWriteEnable,
		input wire csrReadEnable,
		input wire[11:0] csrWriteAddress,
		input wire[11:0] csrReadAddress,
		input wire[31:0] csrWriteData,
		output reg[31:0] csrReadData,
		output wire requestOutput,

		// System interface
		input wire[31:0] programCounter,
		input wire[31:0] currentInstruction,
		input wire[31:0] instruction_memoryAddress,
		input wire[31:0] data_memoryAddress,
		input wire isMachineTimerInterrupt,
		input wire isMachineExternalInterrupt,
		input wire isMachineSoftwareInterrupt,
		input wire isFetchAddressMisaligned,
		input wire isDataAddressMisaligned_load,
		input wire isDataAddressMisaligned_store,
		input wire isJumpMissaligned,
		input wire isFetchAccessFault,
		input wire isDataAccessFault_load,
		input wire isDataAccessFault_store,
		input wire isInvalidInstruction,
		input wire isEBREAK,
		input wire isECALL,
		input wire isFetchAddressBreakpoint,
		input wire isDataAddressBreakpoint,
		input wire[15:0] userInterrupts,
		input wire trapReturn,
		output wire inTrap,
		output wire[31:0] trapVector,
		output wire[31:0] trapReturnVector
	);

	reg machineInterruptEnable;
	reg machinePreviousInterruptEnable;
	wire[31:0] mieValue;
	reg[31:0] mtvecValue;
	reg[31:0] mepcValue;
	reg[31:0] mcauseValue;
	reg[31:0] mtvalValue;
	reg[31:0] mipValue;

	wire[11:0] systemInterrupts = { isMachineExternalInterrupt, 1'b0, 1'b0, 1'b0, 
									isMachineTimerInterrupt, 1'b0, 1'b0, 1'b0, 
									isMachineSoftwareInterrupt, 1'b0, 1'b0, 1'b0 };
	wire[31:0] pendingInterrupts = { userInterrupts, 4'b0000, systemInterrupts } & mieValue;

	wire misalignedInstructionFetch = isFetchAddressMisaligned || isJumpMissaligned;

	reg[30:0] trapCause;
	always @(*) begin
		if (isInterrupt) begin
			case (1'b1)
				isMachineSoftwareInterrupt: trapCause <= 30'd3;
				isMachineTimerInterrupt: trapCause <= 30'd7;
				|userInterrupts: trapCause <= 30'd8;
				isMachineExternalInterrupt: trapCause <= 30'd11;
				default: trapCause <= 30'b0;
			endcase
		end else begin
			case (1'b1)
				isFetchAddressBreakpoint: trapCause <= 30'd3;
				isFetchAccessFault: trapCause <= 30'd1;
				isInvalidInstruction: trapCause <= 30'd2;
				misalignedInstructionFetch: trapCause <= 30'd0;
				isECALL: trapCause <= 30'd11;
				isEBREAK: trapCause <= 30'd3;
				isDataAddressBreakpoint: trapCause <= 30'd3;
				isDataAddressMisaligned_store: trapCause <= 30'd6;
				isDataAddressMisaligned_load: trapCause <= 30'd4;
				isDataAccessFault_store: trapCause <= 30'd7;
				isDataAccessFault_load: trapCause <= 30'd5;				
				default: trapCause <= 30'b0;
			endcase
		end		
	end

	// Misaligned instruction fetch sets trap cause to zero, so needs to be triggered specifically
	wire isException = |trapCause || misalignedInstructionFetch;
	wire isInterrupt = |pendingInterrupts;
	wire isBreakPoint = isEBREAK || isFetchAddressBreakpoint || isDataAddressBreakpoint;
	wire isTrap = isException || isInterrupt;

	assign inTrap = isTrap;

	wire[31:0] mipLoadValue = machineInterruptEnable ? pendingInterrupts : 1'b0;

	reg[31:0] mtvalLoadValue;
	always @(*) begin
		 if (isTrap) begin
			 case (1'b1)
				 isBreakPoint: mtvalLoadValue <= programCounter;
				 isFetchAddressMisaligned: mtvalLoadValue <= instruction_memoryAddress;
				 isDataAddressMisaligned_store || isDataAddressMisaligned_load: mtvalLoadValue <=  data_memoryAddress;
				 isInvalidInstruction: mtvalLoadValue <= currentInstruction;
				 default: mtvalLoadValue <= 32'b0;
			 endcase			
		 end else begin
			 mtvalLoadValue <= 32'b0;
		 end 
	end

	// mstatus
	wire[31:0] mstatusReadData;
	wire mstatusRequestOutput;
	wire mstatusReadDataEnable_nc;
	wire[31:0] mstatusWriteData;
	wire mstatusWriteDataEnable;
	CSR_DataRegister #(.ADDRESS(12'h300)) mstatus(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(mstatusReadData),
		.csrRequestOutput(mstatusRequestOutput),
		.readData( { 25'b0, machinePreviousInterruptEnable, 3'b0, machineInterruptEnable, 2'b0 } ),
		.readDataEnable(mstatusReadDataEnable_nc),
		.writeData(mstatusWriteData),
		.writeDataEnable(mstatusWriteDataEnable));

	always @(posedge clk) begin
		if (rst) begin
			machineInterruptEnable <= 1'b0;
			machinePreviousInterruptEnable <= 1'b0;
		end
		else begin
			if (trapReturn) begin
				machineInterruptEnable <= machinePreviousInterruptEnable;
				machinePreviousInterruptEnable <= 1'b0;
			end else if (isTrap) begin
				machineInterruptEnable <= 1'b0;
				machinePreviousInterruptEnable <= machineInterruptEnable;
			end else if (mstatusWriteDataEnable) begin
				machineInterruptEnable <=  mstatusWriteData[3];
				machinePreviousInterruptEnable <=  mstatusWriteData[7];
			end
		end
	end

	// mie
	wire[31:0] mieReadData;
	wire mieRequestOutput;
	CSR_ConfigurationRegister #(.ADDRESS(12'h304), .DEFAULT(32'b0)) mie(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(mieReadData),
		.csrRequestOutput(mieRequestOutput),
		.value(mieValue));

	// mtvec
	// In theory this is a WARL register, so only legal values can be read,
	// This means that some bits should always be zero, but 
	wire[31:0] mtvecValueValid = mtvecValue;//{ mtvecValue[31:4] , 2'b00, 1'b0, mtvecValue[0] }; 
	wire mtvecRequestOutput;
	wire[31:0] mtvecReadData;
	wire mtvecReadDataEnable_nc;
	wire[31:0] mtvecWriteData;
	wire mtvecWriteDataEnable;
	CSR_DataRegister #(.ADDRESS(12'h305)) mtvec(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(mtvecReadData),
		.csrRequestOutput(mtvecRequestOutput),
		.readData(mtvecValueValid),
		.readDataEnable(mtvecReadDataEnable_nc),
		.writeData(mtvecWriteData),
		.writeDataEnable(mtvecWriteDataEnable));

	always @(posedge clk) begin
		if (rst) mtvecValue <= 32'b0;
		else begin
			if (mtvecWriteDataEnable) mtvecValue <= mtvecWriteData;
		end
	end

	wire[31:0] trapVectorBase = { mtvecValueValid[31:2], 2'b00 };
	wire[1:0] trapVectorMode = mtvecValueValid[1:0];

	assign trapVector = (trapVectorMode == 2'b01) && isInterrupt ? trapVectorBase + {mcauseValue[29:0], 2'b00} : trapVectorBase;

	// mscratch
	wire[31:0] mscratchReadData;
	wire mscratchRequestOutput;
	wire[31:0] mscratchValue_nc;
	CSR_ConfigurationRegister #(.ADDRESS(12'h340), .DEFAULT(32'b0)) mscratch (
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(mscratchReadData),
		.csrRequestOutput(mscratchRequestOutput),
		.value(mscratchValue_nc));

	// mepc
	wire[31:0] mepcReadData;
	wire mepcRequestOutput;
	wire mepcReadDataEnable_nc;
	wire[31:0] mepcWriteData;
	wire mepcWriteDataEnable;
	CSR_DataRegister #(.ADDRESS(12'h341)) mepc(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(mepcReadData),
		.csrRequestOutput(mepcRequestOutput),
		.readData({ mepcValue[31:1], 1'b0 }),
		.readDataEnable(mepcReadDataEnable_nc),
		.writeData(mepcWriteData),
		.writeDataEnable(mepcWriteDataEnable));

	always @(posedge clk) begin
		if (rst) mepcValue <= 32'b0;
		else begin
			if (isTrap) mepcValue <= programCounter;
			else if (mepcWriteDataEnable) mepcValue <= mepcWriteData;
		end
	end

	assign trapReturnVector = mepcValue;

	// mcause
	wire[31:0] mcauseReadData;
	wire mcauseRequestOutput;
	wire mcauseReadDataEnable_nc;
	wire[31:0] mcauseWriteData;
	wire mcauseWriteDataEnable;
	CSR_DataRegister #(.ADDRESS(12'h342)) mcause(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(mcauseReadData),
		.csrRequestOutput(mcauseRequestOutput),
		.readData(mcauseValue),
		.readDataEnable(mcauseReadDataEnable_nc),
		.writeData(mcauseWriteData),
		.writeDataEnable(mcauseWriteDataEnable));

	always @(posedge clk) begin
		if (rst) mcauseValue <= 32'b0;
		else begin
			if (isTrap) mcauseValue <= { isInterrupt, trapCause };
			else if (mcauseWriteDataEnable) mcauseValue <= mcauseWriteData;
		end
	end

	// mtval
	wire[31:0] mtvalReadData;
	wire mtvalRequestOutput;
	wire mtvalReadDataEnable_nc;
	wire[31:0] mtvalWriteData;
	wire mtvalWriteDataEnable;
	CSR_DataRegister #(.ADDRESS(12'h343)) mtval(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(mtvalReadData),
		.csrRequestOutput(mtvalRequestOutput),
		.readData(mtvalValue),
		.readDataEnable(mtvalReadDataEnable_nc),
		.writeData(mtvalWriteData),
		.writeDataEnable(mtvalWriteDataEnable));

	always @(posedge clk) begin
		if (rst) mtvalValue <= 32'b0;
		else begin
			if (isTrap) mtvalValue <= mtvalLoadValue;
			else if (mtvalWriteDataEnable) mtvalValue <= mtvalWriteData;
		end
	end

	// mip
	wire[31:0] mipReadData;
	wire mipRequestOutput;
	wire mipReadDataEnable_nc;
	wire[31:0] mipWriteData;
	wire mipWriteDataEnable;
	CSR_DataRegister #(.ADDRESS(12'h344)) mip(
		.clk(clk),
		.rst(rst),
		.csrWriteEnable(csrWriteEnable),
		.csrReadEnable(csrReadEnable),
		.csrWriteAddress(csrWriteAddress),
		.csrReadAddress(csrReadAddress),
		.csrWriteData(csrWriteData),
		.csrReadData(mipReadData),
		.csrRequestOutput(mipRequestOutput),
		.readData(mipValue),
		.readDataEnable(mipReadDataEnable_nc),
		.writeData(mipWriteData),
		.writeDataEnable(mipWriteDataEnable));

	always @(posedge clk) begin
		if (rst) mipValue <= 32'b0;
		else begin
			if (isTrap && isInterrupt) mipValue <= mipLoadValue;
			else if (mipWriteDataEnable) mipValue <= mipWriteData;
		end
	end

	assign requestOutput = mstatusRequestOutput 
						|| mieRequestOutput 
						|| mtvecRequestOutput 
						|| mscratchRequestOutput 
						|| mepcRequestOutput
						|| mcauseRequestOutput
						|| mtvalRequestOutput
						|| mipRequestOutput;

	always @(*) begin
		case (1'b1)
			mstatusRequestOutput: csrReadData <= mstatusReadData;
			mieRequestOutput: csrReadData <= mieReadData;
			mtvecRequestOutput: csrReadData <= mtvecReadData;
			mscratchRequestOutput: csrReadData <= mscratchReadData;
			mepcRequestOutput: csrReadData <= mepcReadData;
			mcauseRequestOutput: csrReadData <= mcauseReadData;
			mtvalRequestOutput: csrReadData <= mtvalReadData;
			mipRequestOutput: csrReadData <= mipReadData;
			default: csrReadData <= 32'b0;
		endcase
	end

endmodulemodule JTAG (
		input wire clk,
		input wire rst,

		input wire[31:0] coreID,
		input wire[10:0] manufacturerID,
		input wire[15:0] partID,
		input wire[3:0] versionID,

		// JTAG interface
		input wire jtag_tck,
		input wire jtag_tms,
		input wire jtag_tdi,
		output wire jtag_tdo,

		// Management interface
		output wire management_enable,
		output wire management_writeEnable,
		output wire[3:0] management_byteSelect,
		output wire[19:0] management_address,
		output wire[31:0] management_writeData,
		input wire[31:0] management_readData,

		output wire[4:0] probe_jtagInstruction
	);
	
	wire[31:0] idcode = { versionID, partID, manufacturerID, 1'b1 };

	// TAP states
	localparam STATE_TEST_LOGIC_RESET = 4'h0;
	localparam STATE_RUN_TEST_IDLE 	  = 4'h1;
	localparam STATE_DR_SELECT_SCAN   = 4'h2;
	localparam STATE_DR_CAPTURE 	  = 4'h3;
	localparam STATE_DR_SHIFT 		  = 4'h4;
	localparam STATE_DR_EXIT_1 		  = 4'h5;
	localparam STATE_DR_PAUSE 		  = 4'h6;
	localparam STATE_DR_EXIT_2 		  = 4'h7;
	localparam STATE_DR_UPDATE 		  = 4'h8;
	localparam STATE_IR_SELECT_SCAN   = 4'h9;
	localparam STATE_IR_CAPTURE 	  = 4'hA;
	localparam STATE_IR_SHIFT 		  = 4'hB;
	localparam STATE_IR_EXIT_1 		  = 4'hC;
	localparam STATE_IR_PAUSE 		  = 4'hD;
	localparam STATE_IR_EXIT_2 		  = 4'hE;
	localparam STATE_IR_UPDATE 		  = 4'hF;

	// https://www.microsemi.com/document-portal/doc_download/130050-ac160-ieee-standard-1149-1-jtag-in-the-sx-rtsx-sx-a-ex-rt54sx-s-families-app-note
	localparam INSTRUCTION_EXTEST 	= 5'b00000;
	localparam INSTRUCTION_SAMPLE 	= 5'b00001;
	localparam INSTRUCTION_INTEST 	= 5'b00010;
	localparam INSTRUCTION_USERCODE = 5'b00011;
	localparam INSTRUCTION_IDCODE 	= 5'b00100;
	localparam INSTRUCTION_BYPASS 	= 5'b11111;
	
	reg tckState = 1'b0;
	reg tckRisingEdge = 1'b0;
	reg tckFallingEdge = 1'b0;

	always @(posedge clk) begin
		if (rst) begin
			tckState <= 1'b0;
			tckRisingEdge = 1'b0;
			tckFallingEdge = 1'b0;
		end else begin
			if (jtag_tck != tckState) begin
				if (jtag_tck) tckRisingEdge = 1'b1;
				else tckFallingEdge = 1'b1;

				tckState <= jtag_tck;
			end else begin
				tckRisingEdge = 1'b0;
				tckFallingEdge = 1'b0;
			end
		end
	end

	reg[3:0] state = STATE_TEST_LOGIC_RESET;
	wire testReset 	   = state == STATE_TEST_LOGIC_RESET;
	wire irCapture 	   = state == STATE_IR_CAPTURE;
	wire drCapture 	   = state == STATE_DR_CAPTURE;
	wire irShiftEnable = state == STATE_IR_SHIFT;
	wire drShiftEnable = state == STATE_DR_SHIFT;
	wire irUpdate 	   = state == STATE_IR_UPDATE;
	wire drUpdate 	   = state == STATE_DR_UPDATE;

	// Instruction register
	reg[4:0] currentInstruction = INSTRUCTION_IDCODE;
	wire irDataOut;
	wire[4:0] irDataRead;
	JTAGRegister #(.WIDTH(5)) instructionRegister (
		.clk(clk),
		.rst(rst),
		.loadEnable(irCapture && tckRisingEdge),
		.shiftEnable(irShiftEnable && tckRisingEdge),
		.parallelIn(currentInstruction),
		.parallelOut(irDataRead),
		.serialIn(jtag_tdi),
		.serialOut(irDataOut));

	always @(posedge clk) begin
		if (rst) currentInstruction <= INSTRUCTION_IDCODE;
		else if ((irUpdate || testReset) && tckRisingEdge) currentInstruction <= irDataRead;
	end

	// Data registers
	// Boundary scan register
	wire drBSRSelect = currentInstruction == INSTRUCTION_SAMPLE;
	wire bsrReadEnable = drBSRSelect && drCapture && tckRisingEdge;
	wire bsrWriteEnable = drBSRSelect && drUpdate && tckRisingEdge;
	wire drBSRDataOut;
	wire[31:0] bsrDataWrite;
	wire[31:0] bsrDataRead;
	JTAGRegister #(.WIDTH(32)) dataBSRRegister (
		.clk(clk),
		.rst(rst),
		.loadEnable(bsrReadEnable),
		.shiftEnable(drBSRSelect && drShiftEnable && tckRisingEdge),
		.parallelIn(bsrDataWrite),
		.parallelOut(bsrDataRead),
		.serialIn(jtag_tdi),
		.serialOut(drBSRDataOut));

	// Bypass register
	wire drBypassSelect = currentInstruction == INSTRUCTION_BYPASS;
	wire drBypassDataOut;
	wire dataBypassRegisterParallelOut_nc;
	JTAGRegister #(.WIDTH(1)) dataBypassRegister (
		.clk(clk),
		.rst(rst),
		.loadEnable(drBypassSelect && drCapture && tckRisingEdge),
		.shiftEnable(drBypassSelect && drShiftEnable && tckRisingEdge),
		.parallelIn(1'b0),
		.parallelOut(dataBypassRegisterParallelOut_nc),
		.serialIn(jtag_tdi),
		.serialOut(drBypassDataOut));

	// ID code register
	wire drIDUserCode = (currentInstruction == INSTRUCTION_USERCODE);
	wire drIDBaseCode = (currentInstruction == INSTRUCTION_IDCODE);
	wire drIDSelect = drIDUserCode || drIDBaseCode;
	wire[31:0] drIDDataIn = drIDUserCode ? coreID : idcode;
	wire drIDDataOut;
	wire[31:0] dataIDRegisterParallelOut_nc;
	JTAGRegister #(.WIDTH(32)) dataIDRegister (
		.clk(clk),
		.rst(rst),
		.loadEnable(drIDSelect && drCapture && tckRisingEdge),
		.shiftEnable(drIDSelect && drShiftEnable && tckRisingEdge),
		.parallelIn(drIDDataIn),
		.parallelOut(dataIDRegisterParallelOut_nc),
		.serialIn(jtag_tdi),
		.serialOut(drIDDataOut));

	wire drDataOut = drBSRSelect 	? drBSRDataOut : 
					 drBypassSelect ? drBypassDataOut : 
					 drIDSelect 	? drIDDataOut :
					 				  1'b0;

	assign jtag_tdo = drShiftEnable ? drDataOut :
				 	  irShiftEnable ? irDataOut :
				 				 	  1'b0;

	always @(posedge clk) begin
		if (rst) begin
			state <= STATE_TEST_LOGIC_RESET;
		end else begin
			if (tckRisingEdge) begin
				case (state)
					STATE_TEST_LOGIC_RESET:	state <= jtag_tms ? STATE_TEST_LOGIC_RESET : STATE_RUN_TEST_IDLE;
					STATE_RUN_TEST_IDLE:	state <= jtag_tms ? STATE_DR_SELECT_SCAN   : STATE_RUN_TEST_IDLE;
					STATE_DR_SELECT_SCAN:	state <= jtag_tms ? STATE_IR_SELECT_SCAN   : STATE_DR_CAPTURE;
					STATE_DR_CAPTURE:		state <= jtag_tms ? STATE_DR_EXIT_1 	   : STATE_DR_SHIFT;
					STATE_DR_SHIFT:			state <= jtag_tms ? STATE_DR_EXIT_1 	   : STATE_DR_SHIFT;
					STATE_DR_EXIT_1:		state <= jtag_tms ? STATE_DR_UPDATE 	   : STATE_DR_PAUSE;
					STATE_DR_PAUSE:			state <= jtag_tms ? STATE_DR_EXIT_2 	   : STATE_DR_PAUSE;
					STATE_DR_EXIT_2:		state <= jtag_tms ? STATE_DR_UPDATE 	   : STATE_DR_SHIFT;
					STATE_DR_UPDATE:		state <= jtag_tms ? STATE_DR_SELECT_SCAN   : STATE_RUN_TEST_IDLE;
					STATE_IR_SELECT_SCAN:	state <= jtag_tms ? STATE_TEST_LOGIC_RESET : STATE_IR_CAPTURE;
					STATE_IR_CAPTURE:		state <= jtag_tms ? STATE_IR_EXIT_1 	   : STATE_IR_SHIFT;
					STATE_IR_SHIFT:			state <= jtag_tms ? STATE_IR_EXIT_1 	   : STATE_IR_SHIFT;
					STATE_IR_EXIT_1:		state <= jtag_tms ? STATE_IR_UPDATE 	   : STATE_IR_PAUSE;
					STATE_IR_PAUSE:			state <= jtag_tms ? STATE_IR_EXIT_2 	   : STATE_IR_PAUSE;
					STATE_IR_EXIT_2:		state <= jtag_tms ? STATE_IR_UPDATE 	   : STATE_IR_SHIFT;
					STATE_IR_UPDATE:		state <= jtag_tms ? STATE_DR_SELECT_SCAN   : STATE_RUN_TEST_IDLE;
					default:				state <= STATE_TEST_LOGIC_RESET;
				endcase
			end
		end
	end

	assign probe_jtagInstruction = currentInstruction;

	// Core managment control
	localparam MANAGEMENT_STATE_IDLE = 3'h0;
	localparam MANAGEMENT_STATE_READ = 3'h1;
	localparam MANAGEMENT_STATE_RETURN_DATA = 3'h2;
	localparam MANAGEMENT_STATE_GET_DATA = 3'h3;
	localparam MANAGEMENT_STATE_WRITE = 3'h4;

	reg[2:0] managementState = MANAGEMENT_STATE_IDLE;
	reg[31:0] managementReadData = 32'b0;
	reg[25:0] managementAddress = 20'b0;
	reg[31:0] managementWriteData = 32'b0;
	reg[3:0] managementByteSelect = 4'h0;

	wire managementCommandByteSelect = bsrDataRead[29:26];
	wire managementCommandWriteEnable = bsrDataRead[30];
	wire managementCommandReadEnable = bsrDataRead[31];

	always @(posedge clk) begin
		if (rst) begin
			managementState <= MANAGEMENT_STATE_IDLE;
			managementReadData <= 32'b0;
			managementAddress <= 26'b0;
			managementWriteData <= 32'b0;
			managementByteSelect <= 4'h0;
		end else begin
			case (managementState)
				MANAGEMENT_STATE_IDLE: begin
					managementReadData <= 32'b0;
					
					if (bsrWriteEnable) begin
						if (!managementCommandByteSelect) begin
							managementAddress <= bsrDataRead[19:0];
							managementByteSelect <= managementCommandByteSelect;

							if (managementCommandWriteEnable) managementState <= MANAGEMENT_STATE_GET_DATA; 
							if (managementCommandReadEnable) managementState <= MANAGEMENT_STATE_READ;
						end
					end
				end

				MANAGEMENT_STATE_READ: begin
					managementReadData <= management_readData;
					managementState <= MANAGEMENT_STATE_RETURN_DATA;
				end

				MANAGEMENT_STATE_RETURN_DATA: begin
					if (bsrReadEnable) managementState <= MANAGEMENT_STATE_IDLE;
				end

				MANAGEMENT_STATE_GET_DATA: begin
					if (bsrWriteEnable) begin
						managementWriteData <= bsrDataRead;
						managementState <= MANAGEMENT_STATE_WRITE; 
					end
				end

				MANAGEMENT_STATE_WRITE: begin
					managementState <= MANAGEMENT_STATE_IDLE;
				end				

				default: begin
					managementState <= MANAGEMENT_STATE_IDLE;
				end
			endcase
		end
	end

	assign bsrDataWrite = managementReadData;

	assign management_writeEnable = managementState == MANAGEMENT_STATE_WRITE;
	assign management_enable = (managementState == MANAGEMENT_STATE_READ) || (managementState == MANAGEMENT_STATE_WRITE);
	assign management_byteSelect = managementByteSelect;
	assign management_address = managementAddress[19:0];
	assign management_writeData = managementState == MANAGEMENT_STATE_WRITE ? managementReadData : 32'b0;

endmodulemodule JTAGRegister #(
		parameter WIDTH = 8
	)(
		input wire clk,
		input wire rst,

		input wire loadEnable,
		input wire shiftEnable,

		input  wire[WIDTH-1:0] parallelIn,
		output wire[WIDTH-1:0] parallelOut,
		input  wire serialIn,
		output wire serialOut
	);

	reg[WIDTH-1:0] data = {WIDTH{1'b0}};
	wire[WIDTH-1:0] nextData;

	generate
		if (WIDTH == 1) begin
			assign nextData = serialIn;
		end else begin
			assign nextData = { data[WIDTH-2:0], serialIn };
		end
	endgenerate

	always @(posedge clk) begin
		if (rst) data <= {WIDTH{1'b0}};
		else if (loadEnable) data <= parallelIn;
		else if (shiftEnable) data <= nextData;
	end
		
	assign parallelOut = data;
	assign serialOut = data[WIDTH-1];

endmodulemodule LocalMemoryInterface #(
		parameter SRAM_ADDRESS_SIZE = 9
	)(
		input wire clk,
		input wire rst,

		// Core interface
		input wire[23:0] coreAddress,
		input wire[3:0] coreByteSelect,
		input wire coreEnable,
		input wire coreWriteEnable,
		input wire[31:0] coreDataWrite,
		output wire[31:0] coreDataRead,
		output wire coreBusy,

		// WB interface
		input wire[23:0] wbAddress,
		input wire[3:0] wbByteSelect,
		input wire wbEnable,
		input wire wbWriteEnable,
		input wire[31:0] wbDataWrite,
		output wire[31:0] wbDataRead,
		output wire wbBusy,

		// Flash interface
		output wire[22:0] flashAddress,
		output wire[3:0] flashByteSelect,
		output wire flashEnable,
		output wire flashWriteEnable,
		output wire[31:0] flashDataWrite,
		input wire[31:0] flashDataRead,
		input wire flashBusy,

		// SRAM rw port
		output wire clk0, // Port clock
		output wire[1:0] csb0, // active low chip select
		output wire web0, // active low write control
		output wire[3:0] wmask0, // write mask
		output wire[SRAM_ADDRESS_SIZE-1:0] addr0,
		output wire[31:0] din0,
		input  wire[63:0] dout0,

		// SRAM r port
		output wire clk1,
		output wire[1:0] csb1,
		output wire[SRAM_ADDRESS_SIZE-1:0] addr1,
		input  wire[63:0] dout1
	);

	// Core enable pins
	wire coreSRAMEnable = coreAddress[23:SRAM_ADDRESS_SIZE+3] == 'b0 && coreEnable;
	wire coreSRAMWriteEnable = coreSRAMEnable && coreWriteEnable;
	wire coreSRAMReadEnable = coreSRAMEnable && !coreWriteEnable;

	// Wishbone enable pins
	wire wbSRAMEnable = wbAddress[23:SRAM_ADDRESS_SIZE+3] == 'b0 && wbEnable;
	wire wbSRAMWriteEnable = wbSRAMEnable && wbWriteEnable;
	wire wbSRAMReadEnable = wbSRAMEnable && !wbWriteEnable;

	// Generate SRAM control signals
	// Core can always read from read only port
	// Core can always write to read/write port
	// Wishbone can read/write to read/write port, but only if core is not writing to it
	wire[31:0] rwPortReadData;
	wire[31:0] rPortReadData;

	wire rBankSelect;
	wire rwBankSelect;

	// Busy signals
	reg coreReadReady = 1'b0;
	reg lastRBankSelect = 1'b0;
	reg[3:0] lastCoreByteSelect = 4'b0;
	always @(posedge clk) begin
		if (rst) begin
			coreReadReady <= 1'b0;
			lastRBankSelect = 1'b0;
			lastCoreByteSelect = 4'b0;
		end else if (!coreBusy) begin
			coreReadReady <= 1'b0;
			lastRBankSelect = 1'b0;
			lastCoreByteSelect = 4'b0;
		end	else if (coreSRAMReadEnable) begin
			coreReadReady <= 1'b1;
			lastRBankSelect <= rBankSelect;
			lastCoreByteSelect <= coreByteSelect;
		end else begin 
			coreReadReady <= 1'b0;
			lastRBankSelect = 1'b0;
			lastCoreByteSelect <= 4'b0;
		end
	end

	reg wbReadReady = 1'b0;
	reg lastRWBankSelect = 1'b0;
	reg[3:0] lastWBByteSelect = 4'b0;
	always @(posedge clk) begin
		if (rst) begin 
			wbReadReady <= 1'b0;
			lastRWBankSelect <= 1'b0;
			lastWBByteSelect <= 4'b0;
		end else if (wbSRAMReadEnable) begin
			wbReadReady <= 1'b1;
			lastRWBankSelect <= rwBankSelect;
			lastWBByteSelect <= wbByteSelect;
		end else begin
			wbReadReady <= 1'b0;
			lastRWBankSelect <= 1'b0;
			lastWBByteSelect <= 4'b0;
		end
	end

	assign coreBusy = !coreReadReady;
	assign wbBusy = (wbSRAMEnable && coreSRAMWriteEnable) || (wbSRAMReadEnable && !wbReadReady);

	// Read/Write port
	wire rwPortEnable = coreSRAMWriteEnable || wbSRAMWriteEnable || (wbSRAMReadEnable && !wbReadReady);
	wire rwWriteEnable = coreSRAMWriteEnable || (!coreSRAMWriteEnable && wbSRAMWriteEnable);
	wire[SRAM_ADDRESS_SIZE:0] rwAddress = coreSRAMWriteEnable ? coreAddress[SRAM_ADDRESS_SIZE+2:2] :
				   						  wbSRAMEnable        ?   wbAddress[SRAM_ADDRESS_SIZE+2:2] : 'b0;
	assign rwBankSelect = rwAddress[SRAM_ADDRESS_SIZE];

	assign wbDataRead = {
		lastWBByteSelect[3] && wbReadReady ? rwPortReadData[31:24] : ~8'h00,
		lastWBByteSelect[2] && wbReadReady ? rwPortReadData[23:16] : ~8'h00,
		lastWBByteSelect[1] && wbReadReady ? rwPortReadData[15:8]  : ~8'h00,
		lastWBByteSelect[0] && wbReadReady ? rwPortReadData[7:0]   : ~8'h00
	};

	// Read port
	wire rPortEnable = coreSRAMReadEnable && !coreReadReady;
	wire[SRAM_ADDRESS_SIZE:0] rAddress = coreAddress[SRAM_ADDRESS_SIZE+2:2];
	assign rBankSelect = rAddress[SRAM_ADDRESS_SIZE];

	assign coreDataRead = {
		lastCoreByteSelect[3] && coreReadReady ? rPortReadData[31:24] : ~8'h00,
		lastCoreByteSelect[2] && coreReadReady ? rPortReadData[23:16] : ~8'h00,
		lastCoreByteSelect[1] && coreReadReady ? rPortReadData[15:8]  : ~8'h00,
		lastCoreByteSelect[0] && coreReadReady ? rPortReadData[7:0]   : ~8'h00
	};

	// SRAM connections
	assign clk0 = clk;
	assign csb0 = { !(rwPortEnable && rwBankSelect), !(rwPortEnable && !rwBankSelect) };
	assign web0 = !rwWriteEnable;
	assign wmask0 = coreSRAMWriteEnable ? coreByteSelect : 
					wbSRAMWriteEnable   ? wbByteSelect   : 4'b0;
	assign addr0 = rwAddress[SRAM_ADDRESS_SIZE-1:0];
	assign din0 = coreSRAMWriteEnable ? coreDataWrite : 
				  wbSRAMWriteEnable   ? wbDataWrite   : 32'b0;
	assign rwPortReadData = lastRWBankSelect ? dout0[63:32] : dout0[31:0];

	assign clk1 = clk;
	assign csb1 = { !(rPortEnable && rBankSelect), !(rPortEnable && !rBankSelect) };
	assign addr1 = rAddress[SRAM_ADDRESS_SIZE-1:0];
	assign rPortReadData = lastRBankSelect ? dout1[63:32] : dout1[31:0];

endmodulemodule MemoryController (
		input wire clk,
		input wire rst,

		// Instruction cache interface
		input wire[31:0] coreInstructionAddress,
		input wire coreInstructionEnable,
		output reg[31:0] coreInstructionDataRead,
		output reg coreInstructionBusy,

		// Data cache interface
		input wire[31:0] coreDataAddress,
		input wire[3:0] coreDataByteSelect,
		input wire coreDataEnable,
		input wire coreDataWriteEnable,
		input wire[31:0] coreDataDataWrite,
		output reg[31:0] coreDataDataRead,
		output reg coreDataBusy,

		// Local memory interface
		output reg[23:0] localMemoryAddress,
		output reg[3:0] localMemoryByteSelect,
		output reg localMemoryEnable,
		output reg localMemoryWriteEnable,
		output reg[31:0] localMemoryDataWrite,
		input wire[31:0] localMemoryDataRead,
		input wire localMemoryBusy,

		// WB interface
		output reg[27:0] wbAddress,
		output reg[3:0] wbByteSelect,
		output reg wbEnable,
		output reg wbWriteEnable,
		output reg[31:0] wbDataWrite,
		input wire[31:0] wbDataRead,
		input wire wbBusy
	);
	
	localparam LOCAL_MEMORY_ADDRESS = 4'b0000;
	localparam WB_ADDRESS 		    = 4'b0001;

	wire instruction_enableLocalMemory = coreInstructionEnable && (coreInstructionAddress[31:24] == { LOCAL_MEMORY_ADDRESS, 4'b0000 });
	wire data_enableLocalMemory 	   = coreDataEnable && (coreDataAddress[31:24] == { LOCAL_MEMORY_ADDRESS, 4'b0000 });
	wire instruction_enableWB 		   = coreInstructionEnable && (coreInstructionAddress[31:28] == WB_ADDRESS);
	wire data_enableWB 		  		   = coreDataEnable && (coreDataAddress[31:28] == WB_ADDRESS);

	reg last_instruction_enableLocalMemory;
	reg last_data_enableLocalMemory;
	reg last_instruction_enableWB;
	reg last_data_enableWB;

	always @(posedge clk) begin
		if (rst) begin
			last_instruction_enableLocalMemory <= 1'b0;
			last_data_enableLocalMemory <= 1'b0;
			last_instruction_enableWB <= 1'b0;
			last_data_enableWB <= 1'b0;
		end else begin
			last_instruction_enableLocalMemory <= instruction_enableLocalMemory;
			last_data_enableLocalMemory <= data_enableLocalMemory;
			last_instruction_enableWB <= instruction_enableWB;
			last_data_enableWB <= data_enableWB;
		end
	end

	always @(*) begin
		case (1'b1)
			instruction_enableLocalMemory: begin
				localMemoryAddress 	   <= coreInstructionAddress[23:0];
				localMemoryByteSelect  <= 4'b1111;
				localMemoryEnable  	   <= coreInstructionEnable;
				localMemoryWriteEnable <= 1'b0;
				localMemoryDataWrite   <= 32'b0;
			end

			data_enableLocalMemory: begin
				localMemoryAddress 	   <= coreDataAddress[23:0];
				localMemoryByteSelect  <= coreDataByteSelect;
				localMemoryEnable  	   <= coreDataEnable;
				localMemoryWriteEnable <= coreDataWriteEnable;
				localMemoryDataWrite   <= coreDataDataWrite;
			end

			default: begin
				localMemoryAddress 	   <= 24'b0;
				localMemoryByteSelect  <=  4'b0;
				localMemoryEnable  	   <=  1'b0;
				localMemoryWriteEnable <=  1'b0;
				localMemoryDataWrite   <= 32'b0;
			end
		endcase
	end

	always @(*) begin
		case (1'b1)
			instruction_enableWB: begin
				wbAddress 	  <= coreInstructionAddress[27:0];
				wbByteSelect  <= 4'b1111;
				wbEnable  	  <= coreInstructionEnable;
				wbWriteEnable <= 1'b0;
				wbDataWrite   <= 32'b0;
			end

			data_enableWB: begin
				wbAddress 	  <= coreDataAddress[27:0];
				wbByteSelect  <= coreDataByteSelect;
				wbEnable  	  <= coreDataEnable;
				wbWriteEnable <= coreDataWriteEnable;
				wbDataWrite   <= coreDataDataWrite;
			end

			default: begin
				wbAddress 	  <= 28'b0;
				wbByteSelect  <=  4'b0;
				wbEnable  	  <=  1'b0;
				wbWriteEnable <=  1'b0;
				wbDataWrite   <= 32'b0;
			end
		endcase
	end

	always @(*) begin
		case (1'b1)
			last_instruction_enableLocalMemory: begin
				coreInstructionDataRead <= localMemoryDataRead;
				coreInstructionBusy 	<= localMemoryBusy;
			end
			
			last_instruction_enableWB: begin
				coreInstructionDataRead <= wbDataRead;
				coreInstructionBusy 	<= wbBusy;
			end

			default: begin
				coreInstructionDataRead <= ~32'b0;
				coreInstructionBusy 	<= 1'b1;
			end
		endcase
	end

	always @(*) begin
		case (1'b1)
			last_data_enableLocalMemory: begin
				coreDataDataRead <= localMemoryDataRead;
				coreDataBusy 	 <= localMemoryBusy || last_instruction_enableLocalMemory;
			end
			
			last_data_enableWB: begin
				coreDataDataRead <= wbDataRead;
				coreDataBusy  	 <= wbBusy || last_instruction_enableWB;
			end

			default: begin
				coreDataDataRead <= ~32'b0;
				coreDataBusy 	 <= 1'b1;
			end
		endcase
	end

endmodulemodule Core_WBInterface #(
		parameter ADDRESS_WIDTH = 28
	)(
		// Wishbone master interface
		input wire wb_clk_i,
		input wire wb_rst_i,
		output wire wb_cyc_o,
		output wire wb_stb_o,
		output wire wb_we_o,
		output wire[3:0] wb_sel_o,
		output wire[31:0] wb_data_o,
		output wire[ADDRESS_WIDTH-1:0] wb_adr_o,
		input wire wb_ack_i,
		input wire wb_stall_i,
		input wire wb_error_i,
		input wire[31:0] wb_data_i,

		// Memory interface from core
		input wire[ADDRESS_WIDTH-1:0] wbAddress,
		input wire[3:0] wbByteSelect,
		input wire wbEnable,
		input wire wbWriteEnable,
		input wire[31:0] wbDataWrite,
		output wire[31:0] wbDataRead,
		output wire wbBusy
	);

	localparam STATE_IDLE  		  = 2'h0;
	localparam STATE_WRITE_SINGLE = 2'h1;
	localparam STATE_READ_SINGLE  = 2'h2;
	localparam STATE_END 		  = 2'h3;
	
	reg[1:0] state = STATE_IDLE;
	reg[31:0] readDataBuffered;

	reg stb = 1'b0;

	always @(posedge wb_clk_i) begin
		if (wb_rst_i || (wb_error_i && state != STATE_IDLE)) begin
			state <= STATE_IDLE;
			stb <= 1'b0;
			readDataBuffered <= ~32'b0;
		end else begin
			case (state)
				STATE_IDLE: begin
					readDataBuffered <= ~32'b0;

					if (wbEnable) begin
						if (wbWriteEnable) begin
							state <= STATE_WRITE_SINGLE;
							stb <= 1'b1;
						end else begin
							state <= STATE_READ_SINGLE;
							stb <= 1'b1;
						end
					end
				end

				STATE_WRITE_SINGLE: begin
					stb <= 1'b0;
					
					if (wb_ack_i) begin
						state <= STATE_END;
					end
				end

				STATE_READ_SINGLE: begin
					stb <= 1'b0;

					if (wb_ack_i) begin
						state <= STATE_END;
						readDataBuffered <= wb_data_i;
					end
				end

				STATE_END: begin
					state <= STATE_IDLE;
				end
				
				default: begin
					state <= STATE_IDLE;
					stb <= 1'b0;
				end
			endcase
		end
	end

	assign wb_cyc_o = state != STATE_IDLE;
	assign wb_stb_o = stb;

	assign wb_we_o = state == STATE_WRITE_SINGLE;
	assign wb_sel_o = wbByteSelect;
	assign wb_data_o = wbDataWrite;
	assign wb_adr_o = wbAddress;
	
	assign wbDataRead = readDataBuffered;
	assign wbBusy = (state != STATE_IDLE) && (state != STATE_END);

endmodulemodule WB_SRAMInterface (
		input wire[3:0] coreID,

		// Wishbone slave interface to sram
		input wire wb_clk_i,
		input wire wb_rst_i,
		input wire wb_cyc_i,
		input wire wb_stb_i,
		input wire wb_we_i,
		input wire[3:0] wb_sel_i,
		input wire[31:0] wb_data_i,
		input wire[23:0] wb_adr_i,
		output wire wb_ack_o,
		output wire wb_stall_o,
		output wire wb_error_o,
		output wire[31:0] wb_data_o,

		// Memory interface
		output wire[23:0] localMemoryAddress,
		output wire[3:0] localMemoryByteSelect,
		output wire localMemoryEnable,
		output wire localMemoryWriteEnable,
		output wire[31:0] localMemoryDataWrite,
		input wire[31:0] localMemoryDataRead,
		input wire localMemoryBusy,

		// Management interface
		output wire management_enable,
		output wire management_writeEnable,
		output wire[3:0] management_byteSelect,
		output wire[19:0] management_address,
		output wire[31:0] management_writeData,
		input wire[31:0] management_readData,
		input wire management_busy
	);
	
	localparam STATE_IDLE  		  = 2'h0;
	localparam STATE_WRITE_SINGLE = 2'h1;
	localparam STATE_READ_SINGLE  = 2'h2;
	localparam STATE_FINISH 	  = 2'h3;
	
	reg[1:0] state = STATE_IDLE;
	reg[23:0] currentAddress;
	reg[3:0] currentByteSelect;
	reg[31:0] currentDataIn;

	wire isStateReadSingle = state == STATE_READ_SINGLE;
	wire isStateWriteSingle = state == STATE_WRITE_SINGLE;
	wire isStateIdle = state == STATE_IDLE;

	wire[31:0] peripheralBus_dataRead;
	wire peripheralBus_busy;

	reg stall = 1'b0;
	reg acknowledge = 1'b0;
	reg[31:0] dataRead_buffered;
	
	always @(posedge wb_clk_i) begin
		if (wb_rst_i) begin
			state <= STATE_IDLE;
			stall <= 1'b0;
			acknowledge <= 1'b0;
			dataRead_buffered <= ~32'b0;
		end else begin
			case (state)
				STATE_IDLE: begin
					stall <= 1'b0;
					acknowledge <= 1'b0;
					dataRead_buffered <= ~32'b0;

					if (wb_cyc_i) begin
						if (wb_stb_i) begin
							currentAddress <= wb_adr_i;
							currentByteSelect <= wb_sel_i;
							currentDataIn <= wb_data_i;
							stall <= 1'b1;

							if (wb_we_i) begin
								state <= STATE_WRITE_SINGLE;
							end else begin
								state <= STATE_READ_SINGLE;
							end
						end
					end
				end

				STATE_WRITE_SINGLE: begin
					if (!peripheralBus_busy) begin
						state <= STATE_FINISH;
						acknowledge <= 1'b1;
					end
				end

				STATE_READ_SINGLE: begin
					if (!peripheralBus_busy) begin
						state <= STATE_FINISH;
						acknowledge <= 1'b1;
						dataRead_buffered <= peripheralBus_dataRead;
					end
				end

				STATE_FINISH: begin
					state <= STATE_IDLE;
					stall <= 1'b0;
					acknowledge <= 1'b0;
					dataRead_buffered <= ~32'b0;
				end

				default: begin
					state <= STATE_IDLE;
					stall <= 1'b0;
					acknowledge <= 1'b0;
				end
			endcase
		end
	end

	// Connect wishbone bus signals
	assign wb_ack_o = acknowledge;
	assign wb_stall_o = stall;
	assign wb_error_o = 1'b0;

	// Connect to local peripheral bus
	wire peripheralBus_we = isStateWriteSingle;
	wire peripheralBus_oe = isStateReadSingle;
	wire[23:0] peripheralBus_address = !isStateIdle ? currentAddress : 24'b0;
	wire[3:0] peripheralBus_byteSelect = !isStateIdle ? currentByteSelect : 4'b0;
	wire[31:0] peripheralBus_dataWrite = isStateWriteSingle ? wb_data_i : 32'b0;	
	assign wb_data_o = dataRead_buffered;

	// Connect local memory and management interface signals
	assign localMemoryEnable = wb_adr_i[23] == 1'b0 && (peripheralBus_oe || peripheralBus_we);
	assign management_enable = wb_adr_i[23:20] == 4'h8 && (peripheralBus_oe || peripheralBus_we);

	assign localMemoryWriteEnable = localMemoryEnable && peripheralBus_we;
	assign peripheralBus_dataRead = localMemoryEnable ? localMemoryDataRead : 
									management_enable   ? management_readData : ~32'b0;
	assign peripheralBus_busy = (localMemoryEnable && localMemoryBusy) || (management_enable && management_busy);

	assign localMemoryAddress = peripheralBus_address;
	assign localMemoryByteSelect = peripheralBus_byteSelect;
	assign localMemoryDataWrite = peripheralBus_dataWrite;

	assign management_writeEnable = management_enable && peripheralBus_we;
	assign management_address = peripheralBus_address;
	assign management_byteSelect = peripheralBus_byteSelect;
	assign management_writeData = peripheralBus_dataWrite;

endmodulemodule Flash (
	
		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground

		input wire wb_clk_i,
		input wire wb_rst_i,

		// Wishbone interface
		input wire wb_cyc_i,
		input wire wb_stb_i,
		input wire wb_we_i,
		input wire[3:0] wb_sel_i,
		input wire[31:0] wb_data_i,
		input wire[23:0] wb_adr_i,
		output wire wb_ack_o,
		output wire wb_stall_o,
		output wire wb_error_o,
		output wire[31:0] wb_data_o,

		// Flash QSPI
		output wire flash_csb,
		output wire flash_sck,
		output wire flash_io0_we,
		output wire flash_io0_write,
		input wire flash_io0_read,
		output wire flash_io1_we,
		output wire flash_io1_write,
		input wire flash_io1_read,

		// Flash controller SRAM rw port
		output wire sram_clk0,
		output wire sram_csb0,
		output wire sram_web0,
		output wire[3:0] sram_wmask0,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram_addr0,
		output wire[31:0] sram_din0,
		input wire[31:0] sram_dout0,

		// Wishbone SRAM r port
		output wire sram_clk1,
		output wire sram_csb1,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram_addr1,
		input wire[31:0] sram_dout1
	);

	localparam SRAM_ADDRESS_SIZE = 9;

	localparam STATE_STARTUP 	   	 = 2'b00;
	localparam STATE_WRITE_COMMAND 	 = 2'b01;
	localparam STATE_CHANGE_ADDRESS  = 2'b11;
	localparam STATE_READ_CONTINUOUS = 2'b11;
	
	// Wishbone interface
	wire peripheralBus_we;
	wire peripheralBus_oe;
	wire peripheralBus_busy;
	wire[23:0] peripheralBus_address;
	wire[3:0] peripheralBus_byteSelect;
	wire[31:0] peripheralBus_dataRead;
	wire[31:0] peripheralBus_dataWrite;
	WBPeripheralBusInterface wbPeripheralBusInterface(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_stb_i(wb_stb_i),
		.wb_cyc_i(wb_cyc_i),
		.wb_we_i(wb_we_i),
		.wb_sel_i(wb_sel_i),
		.wb_data_i(wb_data_i),
		.wb_adr_i(wb_adr_i),
		.wb_ack_o(wb_ack_o),
		.wb_stall_o(wb_stall_o),
		.wb_error_o(wb_error_o),
		.wb_data_o(wb_data_o),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(peripheralBus_dataRead),
		.peripheralBus_busy(peripheralBus_busy));

	// Flash cache
	wire qspi_enable;
	wire[23:0] qspi_address;
	wire qspi_changeAddress;
	wire qspi_requestData;
	wire[31:0] qspi_readData;
	wire qspi_readDataValid;

	FlashBuffer #(.SRAM_ADDRESS_SIZE(SRAM_ADDRESS_SIZE)) flashBuffer(
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(peripheralBus_dataRead),
		.peripheralBus_busy(peripheralBus_busy),
		.qspi_enable(qspi_enable),
		.qspi_address(qspi_address),
		.qspi_changeAddress(qspi_changeAddress),
		.qspi_requestData(qspi_requestData),
		.qspi_readData(qspi_readData),
		.qspi_readDataValid(qspi_readDataValid),
		.sram_clk0(sram_clk0),
		.sram_csb0(sram_csb0),
		.sram_web0(sram_web0),
		.sram_wmask0(sram_wmask0),
		.sram_addr0(sram_addr0),
		.sram_din0(sram_din0),
		.sram_dout0(sram_dout0),
		.sram_clk1(sram_clk1),
		.sram_csb1(sram_csb1),
		.sram_addr1(sram_addr1),
		.sram_dout1(sram_dout1));

	// QSPI controller
	QSPIDevice qspiDevice (
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.qspi_enable(qspi_enable),
		.qspi_address(qspi_address),
		.qspi_changeAddress(qspi_changeAddress),
		.qspi_requestData(qspi_requestData),
		.qspi_readData(qspi_readData),
		.qspi_readDataValid(qspi_readDataValid),
		.flash_csb(flash_csb),
		.flash_sck(flash_sck),
		.flash_io0_we(flash_io0_we),
		.flash_io0_write(flash_io0_write),
		.flash_io0_read(flash_io0_read),
		.flash_io1_we(flash_io1_we),
		.flash_io1_write(flash_io1_write),
		.flash_io1_read(flash_io1_read));

endmodulemodule FlashBuffer #(
		parameter SRAM_ADDRESS_SIZE = 9
	)(
		input wire clk,
		input wire rst,

		// Peripheral Bus
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		input wire[23:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		input wire[31:0] peripheralBus_dataWrite,
		output reg[31:0] peripheralBus_dataRead,
		output wire peripheralBus_busy,

		// QSPI device
		output wire qspi_enable,
		output wire[23:0] qspi_address,
		output wire qspi_changeAddress,
		output reg qspi_requestData,
		input wire[31:0] qspi_readData,
		input wire qspi_readDataValid,

		// Flash controller SRAM rw port
		output wire sram_clk0,
		output wire sram_csb0,
		output wire sram_web0,
		output wire[3:0] sram_wmask0,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram_addr0,
		output wire[31:0] sram_din0,
		input wire[31:0] sram_dout0,

		// Wishbone SRAM r port
		output wire sram_clk1,
		output wire sram_csb1,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram_addr1,
		input wire[31:0] sram_dout1
	);

	reg[23:0] cachedAddress;
	reg[SRAM_ADDRESS_SIZE:0] cachedCount;
	wire[SRAM_ADDRESS_SIZE:0] nextCachedCount = cachedCount + 1;
	wire[SRAM_ADDRESS_SIZE:0] cachedCountFinal = { 1'b1, {(SRAM_ADDRESS_SIZE){1'b0}} };

	// Select
	wire sramEnable = peripheralBus_address[23:SRAM_ADDRESS_SIZE+2] == {(22-SRAM_ADDRESS_SIZE){1'b0}};
	wire registersEnable = peripheralBus_address[23:12] == 12'h001;
	wire[11:0] localAddress = peripheralBus_address[11:0];

	// Register
	// Configuration register 	Default 0x0
	// b00: enable				Default 0x0
	wire[31:0] configurationRegisterOutputData;
	wire configurationRegisterOutputRequest;
	wire configuration;
	ConfigurationRegister #(.WIDTH(1), .ADDRESS(12'h000), .DEFAULT(1'b0)) configurationRegister(
		.clk(clk),
		.rst(rst),
		.enable(registersEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(configurationRegisterOutputData),
		.requestOutput(configurationRegisterOutputRequest),
		.currentValue(configuration));

	assign qspi_enable = configuration;

	// Base address register 	 Default 0x0
	reg[23:0] baseAddress;
	wire[31:0] baseAddressRegisterOutputData;
	wire baseAddressRegisterOutputRequest;
	wire baseAddressRegisterBusBusy_nc;
	wire[23:0] baseAddressRegisterWriteData;
	wire baseAddressRegisterWriteDataEnable;
	wire baseAddressRegisterReadDataEnable_nc;
	DataRegister #(.WIDTH(24), .ADDRESS(12'h004)) baseAddressRegister(
		.clk(clk),
		.rst(rst),
		.enable(registersEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(baseAddressRegisterBusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(baseAddressRegisterOutputData),
		.requestOutput(baseAddressRegisterOutputRequest),
		.writeData(baseAddressRegisterWriteData),
		.writeData_en(baseAddressRegisterWriteDataEnable),
		.writeData_busy(1'b0),
		.readData(baseAddress),
		.readData_en(baseAddressRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	always @(posedge clk) begin
		if (rst) baseAddress <= 24'b0;
		else if (baseAddressRegisterWriteDataEnable) baseAddress <= baseAddressRegisterWriteData;
	end

	// Cached address register
	wire[31:0] cachedAddressRegisterOutputData;
	wire cachedAddressRegisterOutputRequest;
	wire cachedAddressRegisterBusBusy_nc;
	wire[23:0] cachedAddressRegisterWriteData_nc;
	wire cachedAddressRegisterWriteDataEnable_nc;
	wire cachedAddressRegisterReadDataEnable_nc;
	DataRegister #(.WIDTH(24), .ADDRESS(12'h008)) cachedAddressRegister(
		.clk(clk),
		.rst(rst),
		.enable(registersEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(cachedAddressRegisterBusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(cachedAddressRegisterOutputData),
		.requestOutput(cachedAddressRegisterOutputRequest),
		.writeData(cachedAddressRegisterWriteData_nc),
		.writeData_en(cachedAddressRegisterWriteDataEnable_nc),
		.writeData_busy(1'b0),
		.readData(cachedAddress),
		.readData_en(cachedAddressRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	// Remember that the read data is only valid on the next clock cycle
	reg flashCacheReadReady = 1'b0;
	always @(posedge clk) begin
		if (rst) flashCacheReadReady <= 1'b0;
		else if (peripheralBus_oe && sramEnable) flashCacheReadReady <= 1'b1;
		else flashCacheReadReady <= 1'b0;
	end

	// Assign peripheral read
	always @(*) begin
		case (1'b1)
			configurationRegisterOutputRequest: peripheralBus_dataRead <= configurationRegisterOutputData;
			baseAddressRegisterOutputRequest: peripheralBus_dataRead <= baseAddressRegisterOutputData;
			cachedAddressRegisterOutputRequest: peripheralBus_dataRead <= cachedAddressRegisterOutputData;
			flashCacheReadReady: peripheralBus_dataRead <= sram_dout1;
			default: peripheralBus_dataRead <= 32'b0;
		endcase
	end

	assign peripheralBus_busy = peripheralBus_oe && sramEnable && !flashCacheReadReady;

	// QSPI interface
	always @(posedge clk) begin
		if (rst) begin
			cachedAddress <= 32'b0;
			cachedCount <= {SRAM_ADDRESS_SIZE{1'b0}};
			qspi_requestData <= 1'b0;
		end	else if (baseAddressRegisterWriteDataEnable) begin
			cachedAddress <= { baseAddressRegisterWriteData[23:2], 2'b00 };
			cachedCount <= {SRAM_ADDRESS_SIZE{1'b0}};
			qspi_requestData <= 1'b1;
		end else if (qspi_requestData && qspi_readDataValid) begin
			cachedAddress <= cachedAddress + 4;
			cachedCount <= nextCachedCount;
			qspi_requestData <= nextCachedCount != cachedCountFinal;
		end
	end

	assign qspi_address = baseAddressRegisterWriteData;
	assign qspi_changeAddress = baseAddressRegisterWriteDataEnable;

	// Assign sram port
	// Read/write port
	assign sram_clk0 = clk;
	assign sram_csb0 = !(qspi_requestData && qspi_readDataValid);	// Active low chip enable
	assign sram_web0 = 1'b0;	// Active low write enable (probably keep as always write)
	assign sram_wmask0 = 4'b1111;
	assign sram_addr0 = cachedAddress[SRAM_ADDRESS_SIZE+1:2];
	assign sram_din0 = qspi_readData;

	// Read port
	assign sram_clk1 = clk;
	assign sram_csb1 = !(sramEnable && peripheralBus_oe);
	assign sram_addr1 = peripheralBus_address[SRAM_ADDRESS_SIZE+1:2];

endmodulemodule QSPIDevice (
		input wire clk,
		input wire rst,

		// Cache interface
		input wire qspi_enable,
		input wire[23:0] qspi_address,
		input wire qspi_changeAddress,
		input wire qspi_requestData,
		output wire[31:0] qspi_readData,
		output reg qspi_readDataValid,

		// QSPI interface
		output wire flash_csb,
		output reg flash_sck,
		output wire flash_io0_we,
		output wire flash_io0_write,
		input wire flash_io0_read, 	// Unused
		output wire flash_io1_we,
		output wire flash_io1_write,  // Unused (constant 1'b0)
		input wire flash_io1_read
	);
	
	localparam STATE_IDLE = 2'h0;
	localparam STATE_SETUP = 2'h1;
	localparam STATE_SHIFT = 2'h2;
	localparam STATE_END = 2'h3;

	localparam RESET_NONE = 2'h0;
	localparam RESET_START = 2'h1;
	localparam RESET_WAKE = 2'h2;

	// Assign these as constants to be in a default spi mode
	assign flash_io0_we = 1'b1;
	assign flash_io1_we = 1'b0;
	assign flash_io1_write = 1'b0;

	// State control
	reg[1:0] state = STATE_IDLE;
	wire deviceBusy = state != STATE_IDLE;
	reg[1:0] resetState = RESET_NONE;
	wire resetDevice = resetState != RESET_NONE;
	reg settingAddress = 1'b0;

	reg outputClock = 1'b0;	
	reg[4:0] bitCounter = 5'b0;
	wire[4:0] nextBitCounter = bitCounter + 1;
	
	wire shiftInEnable  = outputClock && deviceBusy;
	wire shiftOutEnable = !outputClock && deviceBusy;

	reg[31:0] registerLoadData;
	wire serialOut;
	wire[31:0] flashData;
	ShiftRegister #(.WIDTH(32)) register (
		.clk(clk),
		.rst(rst),
		.loadEnable((!deviceBusy && qspi_changeAddress) || ((state == STATE_SETUP) && resetDevice)),
		.shiftInEnable(shiftInEnable),
		.shiftOutEnable(shiftOutEnable),
		.msbFirst(1'b1),
		.parallelIn(registerLoadData),
		.parallelOut(flashData),
		.serialIn(flash_io1_read),
		.serialOut(serialOut));

	// Reorder bytes
	assign qspi_readData = { flashData[7:0], flashData[15:8], flashData[23:16], flashData[31:24] };

	always @(*) begin
		case (1'b1)
			resetState == RESET_START: registerLoadData <= { 8'hFF, 8'h00, 8'h00, 8'h00 };
			resetState == RESET_WAKE: registerLoadData <= { 8'hAB, 8'h00, 8'h00, 8'h00 };
			qspi_changeAddress: registerLoadData <= { 8'h03, qspi_address };
			default: registerLoadData <= 32'b0;
		endcase
	end

	always @(posedge clk) begin
		if (rst) begin
			state <= STATE_IDLE;
			outputClock <= 1'b0;
			bitCounter <= 5'b0;
			resetState <= RESET_START;
			settingAddress <= 1'b0;
			qspi_readDataValid <= 1'b0;
		end else begin
			case (state)
				STATE_IDLE: begin
					outputClock <= 1'b0;
					bitCounter <= 5'b0;

					if (qspi_enable) begin
						if (resetDevice || qspi_changeAddress) begin
							state <= STATE_SETUP;
							settingAddress <= qspi_changeAddress;
						end
					end
				end

				STATE_SETUP: begin
					state <= STATE_SHIFT;
					bitCounter <= 5'b0;
					outputClock <= 1'b1;
					qspi_readDataValid <= 1'b0;		
				end

				STATE_SHIFT: begin
					if (!outputClock) begin
						if ((resetDevice && bitCounter == 5'h07) || (bitCounter == 5'h1F)) begin
							state <= STATE_END;
							qspi_readDataValid <= !settingAddress;
						end	else begin
							bitCounter <= nextBitCounter;
							outputClock <= 1'b1;
						end
					end else begin
						outputClock <= 1'b0;
					end

					if (qspi_changeAddress) state <= STATE_IDLE;
				end

				STATE_END: begin
					if (qspi_requestData) state <= STATE_SETUP;
					else state <= STATE_IDLE;

					outputClock <= 1'b0;
					settingAddress <= 1'b0;
					qspi_readDataValid <= 1'b0;
					
					if (resetState == RESET_START) resetState <= RESET_WAKE;
					else resetState <= RESET_NONE;
				end

				default: begin
					state <= STATE_IDLE;
					bitCounter <= 5'b0;
					outputClock <= 1'b0;
					settingAddress <= 1'b0;
					qspi_readDataValid <= 1'b0;
					resetState <= RESET_START;
				end
			endcase
		end
	end

	// Buffer the spi clock by one cycle so that it lines up with when data is sampled
	always @(posedge clk) begin
		if (rst) flash_sck <= 1'b0;
		else flash_sck <= outputClock;
	end

	assign flash_io0_write = serialOut & deviceBusy;
	assign flash_csb = !deviceBusy;

endmodulemodule Peripherals (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		// Wishbone Slave ports
		input wire wb_clk_i,
		input wire wb_rst_i,
		input wire wb_stb_i,
		input wire wb_cyc_i,
		input wire wb_we_i,
		input wire[3:0] wb_sel_i,
		input wire[31:0] wb_data_i,
		input wire[23:0] wb_adr_i,
		output wire wb_ack_o,
		output wire wb_stall_o,
		output wire wb_error_o,
		output wire[31:0] wb_data_o,

		// IOs
		input  wire[(19 + 19)-1:0] io_in,
		output wire[(19 + 19)-1:0] io_out,
		output wire[(19 + 19)-1:0] io_oeb,

		// Caravel UART
		input wire internal_uart_rx,
		output wire internal_uart_tx,

		// JTAG
		output wire jtag_tck,
		output wire jtag_tms,
		output wire jtag_tdi,
		input wire jtag_tdo,

		// Flash
		input wire flash_csb,
		input wire flash_sck,
		input wire flash_io0_we,
		input wire flash_io0_write,
		output wire flash_io0_read,
		input wire flash_io1_we,
		input wire flash_io1_write,
		output wire flash_io1_read,

		// IRQ
		// input wire irq_en,
		// output wire irq_in,
		output wire[9:0] peripheral_irq,

		// VGA
		input wire[1:0] vga_r,
		input wire[1:0] vga_g,
		input wire[1:0] vga_b,
		input wire vga_vsync,
		input wire vga_hsync,

		// Logic Analyzer Signals
		output wire[1:0] probe_blink
	);

	wire irq_en = 1'b0;
	wire irq_in;

	wire peripheralBus_we;
	wire peripheralBus_oe;
	wire peripheralBus_busy;
	wire[23:0] peripheralBus_address;
	wire[3:0] peripheralBus_byteSelect;
	reg[31:0] peripheralBus_dataRead;
	wire[31:0] peripheralBus_dataWrite;

	WBPeripheralBusInterface wbPeripheralBusInterface(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_stb_i(wb_stb_i),
		.wb_cyc_i(wb_cyc_i),
		.wb_we_i(wb_we_i),
		.wb_sel_i(wb_sel_i),
		.wb_data_i(wb_data_i),
		.wb_adr_i(wb_adr_i),
		.wb_ack_o(wb_ack_o),
		.wb_stall_o(wb_stall_o),
		.wb_error_o(wb_error_o),
		.wb_data_o(wb_data_o),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(peripheralBus_busy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(peripheralBus_dataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite));

	wire[31:0] uart_peripheralBus_dataRead;
	wire uart_requestOutput;
	wire[3:0] uart_en;	
	wire[3:0] uart_rx;
	wire[3:0] uart_tx;
	wire[3:0] uart_irq;
	UART #(.ID(8'h00)) uart(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(peripheralBus_busy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(uart_peripheralBus_dataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.requestOutput(uart_requestOutput),
		.uart_en(uart_en),
		.uart_rx(uart_rx),
		.uart_tx(uart_tx),
		.uart_irq(uart_irq));

	assign uart_rx[0] = internal_uart_rx;
	assign internal_uart_tx = uart_tx[0];

	wire[31:0] spi_peripheralBus_dataRead;
	wire spi_requestOutput;
	wire[0:0] spi_en;
	wire[0:0] spi_clk;
	wire[0:0] spi_mosi;
	wire[0:0] spi_miso;
	wire[0:0] spi_cs;
	SPI #(.ID(8'h01)) spi(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(peripheralBus_busy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(spi_peripheralBus_dataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.requestOutput(spi_requestOutput),
		.spi_en(spi_en),
		.spi_clk(spi_clk),
		.spi_mosi(spi_mosi),
		.spi_miso(spi_miso),
		.spi_cs(spi_cs));

	wire[31:0] pwm_peripheralBus_dataRead;
	wire pwm_requestOutput;
	wire[15:0] pwm_en;
	wire[15:0] pwm_out;
	wire[3:0] pwm_irq;
	PWM #(.ID(8'h02)) pwm(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(peripheralBus_busy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(pwm_peripheralBus_dataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.requestOutput(pwm_requestOutput),
		.pwm_en(pwm_en),
		.pwm_out(pwm_out),
		.pwm_irq(pwm_irq));

	wire[31:0] gpio_peripheralBus_dataRead;
	wire gpio_requestOutput;
	wire[(19 + 19)-1:0] gpio_input;
	wire[(19 + 19)-1:0] gpio_output;
	wire[(19 + 19)-1:0] gpio_oe;
	wire[1:0] gpio_irq;
	GPIO #(.ID(8'h03)) gpio(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(peripheralBus_busy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(gpio_peripheralBus_dataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.requestOutput(gpio_requestOutput),
		.gpio_input(gpio_input),
		.gpio_output(gpio_output),
		.gpio_oe(gpio_oe),
		.gpio_irq(gpio_irq));

	IOMultiplexer ioMux(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.uart_en(uart_en[3:1]),
		.uart_rx(uart_rx[3:1]),
		.uart_tx(uart_tx[3:1]),
		.spi_en(spi_en),
		.spi_clk(spi_clk),
		.spi_mosi(spi_mosi),
		.spi_miso(spi_miso),
		.spi_cs(spi_cs),
		.pwm_en(pwm_en[7:0]),
		.pwm_out(pwm_out[7:0]),
		.gpio_input(gpio_input),
		.gpio_output(gpio_output),
		.gpio_oe(gpio_oe),
		.io_in(io_in),
		.io_out(io_out),
		.io_oeb(io_oeb),
		.jtag_tck(jtag_tck),
		.jtag_tms(jtag_tms),
		.jtag_tdi(jtag_tdi),
		.jtag_tdo(jtag_tdo),
		.flash_csb(flash_csb),
		.flash_sck(flash_sck),
		.flash_io0_we(flash_io0_we),
		.flash_io0_write(flash_io0_write),
		.flash_io0_read(flash_io0_read),
		.flash_io1_we(flash_io1_we),
		.flash_io1_write(flash_io1_write),
		.flash_io1_read(flash_io1_read),
		.irq_en(irq_en),
		.irq_in(irq_in),
		.vga_r(vga_r),
		.vga_g(vga_g),
		.vga_b(vga_b),
		.vga_vsync(vga_vsync),
		.vga_hsync(vga_hsync),
		.probe_blink(probe_blink));

	always @(*) begin
		case (1'b1)
			uart_requestOutput: peripheralBus_dataRead <= uart_peripheralBus_dataRead;
			spi_requestOutput:  peripheralBus_dataRead <= spi_peripheralBus_dataRead;
			pwm_requestOutput:  peripheralBus_dataRead <= pwm_peripheralBus_dataRead;
			gpio_requestOutput: peripheralBus_dataRead <= gpio_peripheralBus_dataRead;
			default: 			peripheralBus_dataRead <= ~32'b0;
		endcase
	end

	assign peripheral_irq = { pwm_irq, uart_irq, gpio_irq };

endmodulemodule WBPeripheralBusInterface (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		// Wishbone Slave ports
		input wire wb_clk_i,
		input wire wb_rst_i,
		input wire wb_stb_i,
		input wire wb_cyc_i,
		input wire wb_we_i,
		input wire[3:0] wb_sel_i,
		input wire[31:0] wb_data_i,
		input wire[23:0] wb_adr_i,
		output wire wb_ack_o,
		output wire wb_stall_o,
		output wire wb_error_o,
		output wire[31:0] wb_data_o,

		// Peripheral Bus
		output wire peripheralBus_we,
		output wire peripheralBus_oe,
		input wire peripheralBus_busy,
		output wire[23:0] peripheralBus_address,
		output wire[3:0] peripheralBus_byteSelect,
		input wire[31:0] peripheralBus_dataRead,
		output wire[31:0] peripheralBus_dataWrite
	);
	
	localparam STATE_IDLE  		  = 2'h0;
	localparam STATE_WRITE_SINGLE = 2'h1;
	localparam STATE_READ_SINGLE  = 2'h2;
	localparam STATE_FINISH 	  = 2'h3;
	
	reg[1:0] state = STATE_IDLE;
	reg[23:0] currentAddress;
	reg[3:0] currentByteSelect;
	reg[31:0] currentDataIn;

	reg stall = 1'b0;
	reg acknowledge = 1'b0;
	reg[31:0] dataRead_buffered;

	always @(posedge wb_clk_i) begin
		if (wb_rst_i) begin
			state <= STATE_IDLE;
			stall <= 1'b0;
			acknowledge <= 1'b0;
			dataRead_buffered <= ~32'b0;
		end else begin
			case (state)
				STATE_IDLE: begin
					stall <= 1'b0;
					acknowledge <= 1'b0;
					dataRead_buffered <= ~32'b0;

					if (wb_cyc_i) begin
						if (wb_stb_i) begin
							currentAddress <= wb_adr_i;
							currentByteSelect <= wb_sel_i;
							currentDataIn <= wb_data_i;
							stall <= 1'b1;

							if (wb_we_i) begin
								state <= STATE_WRITE_SINGLE;
							end else begin
								state <= STATE_READ_SINGLE;
							end
						end
					end
				end

				STATE_WRITE_SINGLE: begin
					if (!peripheralBus_busy) begin
						state <= STATE_FINISH;
						acknowledge <= 1'b1;
					end
				end

				STATE_READ_SINGLE: begin
					if (!peripheralBus_busy) begin
						state <= STATE_FINISH;
						acknowledge <= 1'b1;
						dataRead_buffered <= peripheralBus_dataRead;
					end
				end

				STATE_FINISH: begin
					state <= STATE_IDLE;
					stall <= 1'b0;
					acknowledge <= 1'b0;
					dataRead_buffered <= ~32'b0;
				end

				default: begin
					state <= STATE_IDLE;
					stall <= 1'b0;
					acknowledge <= 1'b0;
				end
			endcase
		end
	end

	// Connect wishbone bus signals
	assign wb_ack_o = acknowledge;
	assign wb_stall_o = stall;
	assign wb_error_o = 1'b0;

	// Connect peripheral bus signals
	assign peripheralBus_we = state == STATE_WRITE_SINGLE;
	assign peripheralBus_oe = state == STATE_READ_SINGLE;

	assign peripheralBus_address = state != STATE_IDLE ? currentAddress : 24'b0;
	assign peripheralBus_byteSelect = state != STATE_IDLE ? currentByteSelect : 4'b0;

	assign wb_data_o = dataRead_buffered;
	assign peripheralBus_dataWrite = state == STATE_WRITE_SINGLE ? wb_data_i : 32'b0;

endmodulemodule GPIO #(
		parameter ID = 8'h03
	)(

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		input wire clk,
		input wire rst,
		
		// Peripheral Bus
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[23:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,

		input wire[(19 + 19)-1:0] gpio_input,
		output wire[(19 + 19)-1:0] gpio_output,
		output wire[(19 + 19)-1:0] gpio_oe,
		output wire[1:0] gpio_irq
	);
	
	wire[19-1:0] gpio0_input;
	wire[19-1:0] gpio0_output;
	wire[19-1:0] gpio0_oe;
	wire[19-1:0] gpio1_input;
	wire[19-1:0] gpio1_output;
	wire[19-1:0] gpio1_oe;

	// Peripheral select
	wire[15:0] localAddress;
	wire peripheralEnable;
	PeripheralSelect #(.ID(ID)) select(
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.peripheralEnable(peripheralEnable));

	wire[31:0] device0OutputData;
	wire device0OutputRequest;
	wire device0BusBusy_nc;
	GPIODevice #(.ID(4'h1), .IO_COUNT(19)) device0(
		.clk(clk),
		.rst(rst),
		.peripheralEnable(peripheralEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(device0BusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(device0OutputData),
		.requestOutput(device0OutputRequest),
		.gpio_input(gpio0_input),
		.gpio_output(gpio0_output),
		.gpio_oe(gpio0_oe),
		.gpio_irq(gpio_irq[0]));

	wire[31:0] device1OutputData;
	wire device1OutputRequest;
	wire device1BusBusy_nc;
	GPIODevice #(.ID(4'h2), .IO_COUNT(19)) device1(
		.clk(clk),
		.rst(rst),
		.peripheralEnable(peripheralEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(device1BusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(device1OutputData),
		.requestOutput(device1OutputRequest),
		.gpio_input(gpio1_input),
		.gpio_output(gpio1_output),
		.gpio_oe(gpio1_oe),
		.gpio_irq(gpio_irq[1]));

	assign requestOutput = device0OutputRequest || device1OutputRequest;
	assign peripheralBus_dataRead = device0OutputRequest ? device0OutputData :
								    device1OutputRequest ? device1OutputData :
													       ~32'b0;
	assign peripheralBus_busy = 1'b0;

	assign gpio0_input = gpio_input[19-1:0];
	assign gpio1_input = gpio_input[(19 + 19)-1:19];
	assign gpio_output = { gpio1_output, gpio0_output };
	assign gpio_oe = { gpio1_oe, gpio0_oe };

endmodulemodule GPIODevice #(
		parameter ID = 4'h0,
		parameter IO_COUNT = 16
	)(
		input wire clk,
		input wire rst,

		// Peripheral bus
		input wire peripheralEnable,
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[15:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,
		
		// GPIO
		input wire[IO_COUNT-1:0] gpio_input,
		output wire[IO_COUNT-1:0] gpio_output,
		output wire[IO_COUNT-1:0] gpio_oe,
		output reg gpio_irq
	);

	reg[IO_COUNT-1:0] inputBuffered;
	always @(posedge clk) begin
		if (rst) inputBuffered <= {IO_COUNT{1'b0}};
		else inputBuffered <= gpio_input;
	end

	// Device select
	wire[11:0] localAddress;
	wire deviceEnable;
	DeviceSelect #(.ID(ID)) select(
		.peripheralEnable(peripheralEnable),
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.deviceEnable(deviceEnable));

	// Registers
	// OE register: Default 0x0
	wire[31:0] oeRegisterOutputData;
	wire oeRegisterOutputRequest;
	OutputRegister #(.WIDTH(IO_COUNT), .ADDRESS(8'h00), .DEFAULT(~{IO_COUNT{1'b0}})) oeRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(oeRegisterOutputData),
		.requestOutput(oeRegisterOutputRequest),
		.currentValue(gpio_oe));

	// Output data register: Default 0x0
	wire[31:0] outputRegisterOutputData;
	wire outputRegisterOutputRequest;
	OutputRegister #(.WIDTH(IO_COUNT), .ADDRESS(8'h01), .DEFAULT({IO_COUNT{1'b0}})) outputRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(outputRegisterOutputData),
		.requestOutput(outputRegisterOutputRequest),
		.currentValue(gpio_output));

	// Input data register
	wire[31:0] inputRegisterOutputData;
	wire inputRegisterOutputRequest;
	wire inputRegisterBusBusy_nc;
	wire[IO_COUNT-1:0] inputRegisterWriteData_nc;
	wire inputRegisterWriteDataEnable_nc;
	wire inputRegisterReadDataEnable_nc;
	DataRegister #(.WIDTH(IO_COUNT), .ADDRESS(12'h020)) inputRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(inputRegisterBusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(inputRegisterOutputData),
		.requestOutput(inputRegisterOutputRequest),
		.writeData(inputRegisterWriteData_nc),
		.writeData_en(inputRegisterWriteDataEnable_nc),
		.writeData_busy(1'b0),
		.readData(inputBuffered),
		.readData_en(inputRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	// IRQ register: Default 0x0
	wire[31:0] irqEnableRegisterOutputData;
	wire irqEnableRegisterOutputRequest;
	wire[IO_COUNT-1:0] irqEnable;
	OutputRegister #(.WIDTH(IO_COUNT), .ADDRESS(8'h03), .DEFAULT({IO_COUNT{1'b0}})) irqEnableRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(irqEnableRegisterOutputData),
		.requestOutput(irqEnableRegisterOutputRequest),
		.currentValue(irqEnable));

	assign requestOutput = oeRegisterOutputRequest || outputRegisterOutputRequest || inputRegisterOutputRequest || irqEnableRegisterOutputRequest;
	assign peripheralBus_dataRead = oeRegisterOutputRequest 	   ? oeRegisterOutputData :
								    outputRegisterOutputRequest    ? outputRegisterOutputData :
								    inputRegisterOutputRequest     ? inputRegisterOutputData :
									irqEnableRegisterOutputRequest ? irqEnableRegisterOutputData :
								   								     ~32'b0;
	assign peripheralBus_busy = 1'b0;
	

	wire[IO_COUNT-1:0] pinIRQ = irqEnable & gpio_oe & inputBuffered;

	always @(posedge clk) begin
		if (rst) gpio_irq <= 1'b0;
		else gpio_irq <= |pinIRQ;
	end

endmodulemodule IOMultiplexer (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		input wire clk,
		input wire rst,

		// IO Modules
		// UART
		input wire[3:1] uart_en,
		output wire[3:1] uart_rx,
		input  wire[3:1] uart_tx,

		// SPI
		input wire[0:0] spi_en,
		input wire[0:0] spi_clk,
		input wire[0:0] spi_mosi,
		output wire[0:0] spi_miso,
		input  wire[0:0] spi_cs,

		// PWM
		input wire[7:0] pwm_en,
		input wire[7:0] pwm_out,

		// GPIO
		output wire[(19 + 19)-1:0] gpio_input,
		input  wire[(19 + 19)-1:0] gpio_output,
		input  wire[(19 + 19)-1:0] gpio_oe,

		// IO Pads
    	input  wire[(19 + 19)-1:0] io_in,
    	output wire[(19 + 19)-1:0] io_out,
    	output wire[(19 + 19)-1:0] io_oeb,

		// JTAG
		output wire jtag_tck,
		output wire jtag_tms,
		output wire jtag_tdi,
		input wire jtag_tdo,

		// Flash
		input wire flash_csb,
		input wire flash_sck,
		input wire flash_io0_we,
		input wire flash_io0_write,
		output wire flash_io0_read,
		input wire flash_io1_we,
		input wire flash_io1_write,
		output wire flash_io1_read,

		// IRQ
		input wire irq_en,
		output wire irq_in,

		// VGA
		input wire[1:0] vga_r,
		input wire[1:0] vga_g,
		input wire[1:0] vga_b,
		input wire vga_vsync,
		input wire vga_hsync,

		output wire[1:0] probe_blink
	);

	// Test blink
	localparam BLINK_CLOCK_DIV = 26;
	reg blinkEnabled = 1'b1;
	wire[1:0] blink;
	Counter #(.WIDTH(2), .DIV(BLINK_CLOCK_DIV), .TOP(0)) ctr(.clk(clk), .rst(rst), .halt(1'b0), .value(blink));

	always @(posedge clk) begin
		if (rst) blinkEnabled <= 1'b1;
		else if (gpio_oe[PIN_BLINK0]) blinkEnabled <= 1'b0;
	end

	assign probe_blink = blink;

	wire jtag;
	wire sdo;
	wire sdi;
	wire csb;
	wire sck;

	assign jtag_tck = sck;
	assign jtag_tms = csb;
	assign jtag_tdi = sdi;
	assign sdo = jtag_tdo;

	//-------------------------------------------------//
	//----------------Pin Mapping Start----------------//
	//-------------Start of Generated Code-------------//

	// Interface IO mapping
	// GPIO0 (user1 side)
	// IO00: JTAG
	// IO01: SDO
	// IO02: SDI
	// IO03: CSB
	// IO04: SCK
	// IO05: GPIO05 or UART1_RX
	// IO06: GPIO06 or UART1_TX
	// IO07: GPIO07 or IRQ
	// IO08: FLASH_CSB
	// IO09: FLASH_SCK
	// IO10: FLASH_IO0
	// IO11: FLASH_IO1
	// IO12: GPIO12 or PWM0
	// IO13: GPIO13 or PWM1
	// IO14: GPIO14 or PWM2
	// IO15: GPIO15 or PWM3
	// IO16: GPIO16 or PWM4
	// IO17: GPIO17 or PWM5
	// IO18: GPIO18 or PWM6

	// GPIO1 (user2 side)
	// IO19: GPIO19 or UART2_RX
	// IO20: GPIO20 or UART2_TX
	// IO21: GPIO21 or PWM7
	// IO22: GPIO22 or SPI0_CLK
	// IO23: GPIO23 or SPI0_MOSI
	// IO24: GPIO24 or SPI0_MISO
	// IO25: GPIO25 or SPI0_CS
	// IO26: GPIO26 or UART3_RX
	// IO27: GPIO27 or UART3_TX
	// IO28: GPIO28 or BLINK0
	// IO29: GPIO29 or BLINK1
	// IO30: VGA_R0
	// IO31: VGA_R1
	// IO32: VGA_G0
	// IO33: VGA_G1
	// IO34: VGA_B0
	// IO35: VGA_B1
	// IO36: VGA_VSYNC
	// IO37: VGA_HSYNC
	
	// IO00-PIN_JTAG: Input
	localparam PIN_JTAG = 0;
	assign gpio_input[PIN_JTAG] = 1'b0;
	assign io_out[PIN_JTAG] = 1'b0;
	assign io_oeb[PIN_JTAG] = 1'b1;
	assign jtag = io_in[PIN_JTAG];
	
	// IO01-PIN_SDO: Output
	localparam PIN_SDO = 1;
	assign gpio_input[PIN_SDO] = 1'b0;
	assign io_out[PIN_SDO] = sdo;
	assign io_oeb[PIN_SDO] = 1'b0;
	
	// IO02-PIN_SDI: Input
	localparam PIN_SDI = 2;
	assign gpio_input[PIN_SDI] = 1'b0;
	assign io_out[PIN_SDI] = 1'b0;
	assign io_oeb[PIN_SDI] = 1'b1;
	assign sdi = io_in[PIN_SDI];
	
	// IO03-PIN_CSB: Input
	localparam PIN_CSB = 3;
	assign gpio_input[PIN_CSB] = 1'b0;
	assign io_out[PIN_CSB] = 1'b0;
	assign io_oeb[PIN_CSB] = 1'b1;
	assign csb = io_in[PIN_CSB];
	
	// IO04-PIN_SCK: Input
	localparam PIN_SCK = 4;
	assign gpio_input[PIN_SCK] = 1'b0;
	assign io_out[PIN_SCK] = 1'b0;
	assign io_oeb[PIN_SCK] = 1'b1;
	assign sck = io_in[PIN_SCK];
	
	// IO05-PIN_UART1_RX: Input
	localparam PIN_UART1_RX = 5;
	assign gpio_input[PIN_UART1_RX] = uart_en[1] ? 1'b0 : (gpio_oe[PIN_UART1_RX] ? io_in[PIN_UART1_RX] : 1'b0);
	assign io_out[PIN_UART1_RX] = uart_en[1] ? 1'b0 : gpio_output[PIN_UART1_RX];
	assign io_oeb[PIN_UART1_RX] = uart_en[1] ? 1'b1 : gpio_oe[PIN_UART1_RX];
	assign uart_rx[1] = uart_en[1] ? io_in[PIN_UART1_RX] : 1'b1;
	
	// IO06-PIN_UART1_TX: Output
	localparam PIN_UART1_TX = 6;
	assign gpio_input[PIN_UART1_TX] = uart_en[1] ? 1'b0 : (gpio_oe[PIN_UART1_TX] ? io_in[PIN_UART1_TX] : 1'b0);
	assign io_out[PIN_UART1_TX] = uart_en[1] ? uart_tx[1] : gpio_output[PIN_UART1_TX];
	assign io_oeb[PIN_UART1_TX] = uart_en[1] ? 1'b0 : gpio_oe[PIN_UART1_TX];
	
	// IO07-PIN_IRQ: Input
	localparam PIN_IRQ = 7;
	assign gpio_input[PIN_IRQ] = irq_en ? 1'b0 : (gpio_oe[PIN_IRQ] ? io_in[PIN_IRQ] : 1'b0);
	assign io_out[PIN_IRQ] = irq_en ? 1'b0 : gpio_output[PIN_IRQ];
	assign io_oeb[PIN_IRQ] = irq_en ? 1'b1 : gpio_oe[PIN_IRQ];
	assign irq_in = irq_en ? io_in[PIN_IRQ] : 1'b0;
	
	// IO08-PIN_FLASH_CSB: Output
	localparam PIN_FLASH_CSB = 8;
	assign gpio_input[PIN_FLASH_CSB] = 1'b0;
	assign io_out[PIN_FLASH_CSB] = flash_csb;
	assign io_oeb[PIN_FLASH_CSB] = 1'b0;
	
	// IO09-PIN_FLASH_SCK: Output
	localparam PIN_FLASH_SCK = 9;
	assign gpio_input[PIN_FLASH_SCK] = 1'b0;
	assign io_out[PIN_FLASH_SCK] = flash_sck;
	assign io_oeb[PIN_FLASH_SCK] = 1'b0;
	
	// IO10-PIN_FLASH_IO0: InOut
	localparam PIN_FLASH_IO0 = 10;
	assign gpio_input[PIN_FLASH_IO0] = 1'b0;
	assign io_out[PIN_FLASH_IO0] = flash_io0_write;
	assign io_oeb[PIN_FLASH_IO0] = !flash_io0_we;
	assign flash_io0_read = !flash_io0_we ? io_in[PIN_FLASH_IO0] : 1'b0;
	
	// IO11-PIN_FLASH_IO1: InOut
	localparam PIN_FLASH_IO1 = 11;
	assign gpio_input[PIN_FLASH_IO1] = 1'b0;
	assign io_out[PIN_FLASH_IO1] = flash_io1_write;
	assign io_oeb[PIN_FLASH_IO1] = !flash_io1_we;
	assign flash_io1_read = !flash_io1_we ? io_in[PIN_FLASH_IO1] : 1'b0;
	
	// IO12-PIN_PWM0: Output
	localparam PIN_PWM0 = 12;
	assign gpio_input[PIN_PWM0] = pwm_en[0] ? 1'b0 : (gpio_oe[PIN_PWM0] ? io_in[PIN_PWM0] : 1'b0);
	assign io_out[PIN_PWM0] = pwm_en[0] ? pwm_out[0] : gpio_output[PIN_PWM0];
	assign io_oeb[PIN_PWM0] = pwm_en[0] ? 1'b0 : gpio_oe[PIN_PWM0];
	
	// IO13-PIN_PWM1: Output
	localparam PIN_PWM1 = 13;
	assign gpio_input[PIN_PWM1] = pwm_en[1] ? 1'b0 : (gpio_oe[PIN_PWM1] ? io_in[PIN_PWM1] : 1'b0);
	assign io_out[PIN_PWM1] = pwm_en[1] ? pwm_out[1] : gpio_output[PIN_PWM1];
	assign io_oeb[PIN_PWM1] = pwm_en[1] ? 1'b0 : gpio_oe[PIN_PWM1];
	
	// IO14-PIN_PWM2: Output
	localparam PIN_PWM2 = 14;
	assign gpio_input[PIN_PWM2] = pwm_en[2] ? 1'b0 : (gpio_oe[PIN_PWM2] ? io_in[PIN_PWM2] : 1'b0);
	assign io_out[PIN_PWM2] = pwm_en[2] ? pwm_out[2] : gpio_output[PIN_PWM2];
	assign io_oeb[PIN_PWM2] = pwm_en[2] ? 1'b0 : gpio_oe[PIN_PWM2];
	
	// IO15-PIN_PWM3: Output
	localparam PIN_PWM3 = 15;
	assign gpio_input[PIN_PWM3] = pwm_en[3] ? 1'b0 : (gpio_oe[PIN_PWM3] ? io_in[PIN_PWM3] : 1'b0);
	assign io_out[PIN_PWM3] = pwm_en[3] ? pwm_out[3] : gpio_output[PIN_PWM3];
	assign io_oeb[PIN_PWM3] = pwm_en[3] ? 1'b0 : gpio_oe[PIN_PWM3];
	
	// IO16-PIN_PWM4: Output
	localparam PIN_PWM4 = 16;
	assign gpio_input[PIN_PWM4] = pwm_en[4] ? 1'b0 : (gpio_oe[PIN_PWM4] ? io_in[PIN_PWM4] : 1'b0);
	assign io_out[PIN_PWM4] = pwm_en[4] ? pwm_out[4] : gpio_output[PIN_PWM4];
	assign io_oeb[PIN_PWM4] = pwm_en[4] ? 1'b0 : gpio_oe[PIN_PWM4];
	
	// IO17-PIN_PWM5: Output
	localparam PIN_PWM5 = 17;
	assign gpio_input[PIN_PWM5] = pwm_en[5] ? 1'b0 : (gpio_oe[PIN_PWM5] ? io_in[PIN_PWM5] : 1'b0);
	assign io_out[PIN_PWM5] = pwm_en[5] ? pwm_out[5] : gpio_output[PIN_PWM5];
	assign io_oeb[PIN_PWM5] = pwm_en[5] ? 1'b0 : gpio_oe[PIN_PWM5];
	
	// IO18-PIN_PWM6: Output
	localparam PIN_PWM6 = 18;
	assign gpio_input[PIN_PWM6] = pwm_en[6] ? 1'b0 : (gpio_oe[PIN_PWM6] ? io_in[PIN_PWM6] : 1'b0);
	assign io_out[PIN_PWM6] = pwm_en[6] ? pwm_out[6] : gpio_output[PIN_PWM6];
	assign io_oeb[PIN_PWM6] = pwm_en[6] ? 1'b0 : gpio_oe[PIN_PWM6];
	
	// IO19-PIN_UART2_RX: Input
	localparam PIN_UART2_RX = 19;
	assign gpio_input[PIN_UART2_RX] = uart_en[2] ? 1'b0 : (gpio_oe[PIN_UART2_RX] ? io_in[PIN_UART2_RX] : 1'b0);
	assign io_out[PIN_UART2_RX] = uart_en[2] ? 1'b0 : gpio_output[PIN_UART2_RX];
	assign io_oeb[PIN_UART2_RX] = uart_en[2] ? 1'b1 : gpio_oe[PIN_UART2_RX];
	assign uart_rx[2] = uart_en[2] ? io_in[PIN_UART2_RX] : 1'b1;
	
	// IO20-PIN_UART2_TX: Output
	localparam PIN_UART2_TX = 20;
	assign gpio_input[PIN_UART2_TX] = uart_en[2] ? 1'b0 : (gpio_oe[PIN_UART2_TX] ? io_in[PIN_UART2_TX] : 1'b0);
	assign io_out[PIN_UART2_TX] = uart_en[2] ? uart_tx[2] : gpio_output[PIN_UART2_TX];
	assign io_oeb[PIN_UART2_TX] = uart_en[2] ? 1'b0 : gpio_oe[PIN_UART2_TX];
	
	// IO21-PIN_PWM7: Output
	localparam PIN_PWM7 = 21;
	assign gpio_input[PIN_PWM7] = pwm_en[7] ? 1'b0 : (gpio_oe[PIN_PWM7] ? io_in[PIN_PWM7] : 1'b0);
	assign io_out[PIN_PWM7] = pwm_en[7] ? pwm_out[7] : gpio_output[PIN_PWM7];
	assign io_oeb[PIN_PWM7] = pwm_en[7] ? 1'b0 : gpio_oe[PIN_PWM7];
	
	// IO22-PIN_SPI0_CLK: Output
	localparam PIN_SPI0_CLK = 22;
	assign gpio_input[PIN_SPI0_CLK] = spi_en[0] ? 1'b0 : (gpio_oe[PIN_SPI0_CLK] ? io_in[PIN_SPI0_CLK] : 1'b0);
	assign io_out[PIN_SPI0_CLK] = spi_en[0] ? spi_clk[0] : gpio_output[PIN_SPI0_CLK];
	assign io_oeb[PIN_SPI0_CLK] = spi_en[0] ? 1'b0 : gpio_oe[PIN_SPI0_CLK];
	
	// IO23-PIN_SPI0_MOSI: Output
	localparam PIN_SPI0_MOSI = 23;
	assign gpio_input[PIN_SPI0_MOSI] = spi_en[0] ? 1'b0 : (gpio_oe[PIN_SPI0_MOSI] ? io_in[PIN_SPI0_MOSI] : 1'b0);
	assign io_out[PIN_SPI0_MOSI] = spi_en[0] ? spi_mosi[0] : gpio_output[PIN_SPI0_MOSI];
	assign io_oeb[PIN_SPI0_MOSI] = spi_en[0] ? 1'b0 : gpio_oe[PIN_SPI0_MOSI];
	
	// IO24-PIN_SPI0_MISO: Input
	localparam PIN_SPI0_MISO = 24;
	assign gpio_input[PIN_SPI0_MISO] = spi_en[0] ? 1'b0 : (gpio_oe[PIN_SPI0_MISO] ? io_in[PIN_SPI0_MISO] : 1'b0);
	assign io_out[PIN_SPI0_MISO] = spi_en[0] ? 1'b0 : gpio_output[PIN_SPI0_MISO];
	assign io_oeb[PIN_SPI0_MISO] = spi_en[0] ? 1'b1 : gpio_oe[PIN_SPI0_MISO];
	assign spi_miso[0] = spi_en[0] ? io_in[PIN_SPI0_MISO] : 1'b0;
	
	// IO25-PIN_SPI0_CS: Output
	localparam PIN_SPI0_CS = 25;
	assign gpio_input[PIN_SPI0_CS] = spi_en[0] ? 1'b0 : (gpio_oe[PIN_SPI0_CS] ? io_in[PIN_SPI0_CS] : 1'b0);
	assign io_out[PIN_SPI0_CS] = spi_en[0] ? spi_cs[0] : gpio_output[PIN_SPI0_CS];
	assign io_oeb[PIN_SPI0_CS] = spi_en[0] ? 1'b0 : gpio_oe[PIN_SPI0_CS];
	
	// IO26-PIN_UART3_RX: Input
	localparam PIN_UART3_RX = 26;
	assign gpio_input[PIN_UART3_RX] = uart_en[3] ? 1'b0 : (gpio_oe[PIN_UART3_RX] ? io_in[PIN_UART3_RX] : 1'b0);
	assign io_out[PIN_UART3_RX] = uart_en[3] ? 1'b0 : gpio_output[PIN_UART3_RX];
	assign io_oeb[PIN_UART3_RX] = uart_en[3] ? 1'b1 : gpio_oe[PIN_UART3_RX];
	assign uart_rx[3] = uart_en[3] ? io_in[PIN_UART3_RX] : 1'b1;
	
	// IO27-PIN_UART3_TX: Output
	localparam PIN_UART3_TX = 27;
	assign gpio_input[PIN_UART3_TX] = uart_en[3] ? 1'b0 : (gpio_oe[PIN_UART3_TX] ? io_in[PIN_UART3_TX] : 1'b0);
	assign io_out[PIN_UART3_TX] = uart_en[3] ? uart_tx[3] : gpio_output[PIN_UART3_TX];
	assign io_oeb[PIN_UART3_TX] = uart_en[3] ? 1'b0 : gpio_oe[PIN_UART3_TX];
	
	// IO28-PIN_BLINK0: Output
	localparam PIN_BLINK0 = 28;
	assign gpio_input[PIN_BLINK0] = blinkEnabled ? 1'b0 : (gpio_oe[PIN_BLINK0] ? io_in[PIN_BLINK0] : 1'b0);
	assign io_out[PIN_BLINK0] = blinkEnabled ? blink[0] : gpio_output[PIN_BLINK0];
	assign io_oeb[PIN_BLINK0] = blinkEnabled ? 1'b0 : gpio_oe[PIN_BLINK0];
	
	// IO29-PIN_BLINK1: Output
	localparam PIN_BLINK1 = 29;
	assign gpio_input[PIN_BLINK1] = blinkEnabled ? 1'b0 : (gpio_oe[PIN_BLINK1] ? io_in[PIN_BLINK1] : 1'b0);
	assign io_out[PIN_BLINK1] = blinkEnabled ? blink[1] : gpio_output[PIN_BLINK1];
	assign io_oeb[PIN_BLINK1] = blinkEnabled ? 1'b0 : gpio_oe[PIN_BLINK1];
	
	// IO30-PIN_VGA_R0: Output
	localparam PIN_VGA_R0 = 30;
	assign gpio_input[PIN_VGA_R0] = 1'b0;
	assign io_out[PIN_VGA_R0] = vga_r[0];
	assign io_oeb[PIN_VGA_R0] = 1'b0;
	
	// IO31-PIN_VGA_R1: Output
	localparam PIN_VGA_R1 = 31;
	assign gpio_input[PIN_VGA_R1] = 1'b0;
	assign io_out[PIN_VGA_R1] = vga_r[1];
	assign io_oeb[PIN_VGA_R1] = 1'b0;
	
	// IO32-PIN_VGA_G0: Output
	localparam PIN_VGA_G0 = 32;
	assign gpio_input[PIN_VGA_G0] = 1'b0;
	assign io_out[PIN_VGA_G0] = vga_g[0];
	assign io_oeb[PIN_VGA_G0] = 1'b0;
	
	// IO33-PIN_VGA_G1: Output
	localparam PIN_VGA_G1 = 33;
	assign gpio_input[PIN_VGA_G1] = 1'b0;
	assign io_out[PIN_VGA_G1] = vga_g[1];
	assign io_oeb[PIN_VGA_G1] = 1'b0;
	
	// IO34-PIN_VGA_B0: Output
	localparam PIN_VGA_B0 = 34;
	assign gpio_input[PIN_VGA_B0] = 1'b0;
	assign io_out[PIN_VGA_B0] = vga_b[0];
	assign io_oeb[PIN_VGA_B0] = 1'b0;
	
	// IO35-PIN_VGA_B1: Output
	localparam PIN_VGA_B1 = 35;
	assign gpio_input[PIN_VGA_B1] = 1'b0;
	assign io_out[PIN_VGA_B1] = vga_b[1];
	assign io_oeb[PIN_VGA_B1] = 1'b0;
	
	// IO36-PIN_VGA_VSYNC: Output
	localparam PIN_VGA_VSYNC = 36;
	assign gpio_input[PIN_VGA_VSYNC] = 1'b0;
	assign io_out[PIN_VGA_VSYNC] = vga_vsync;
	assign io_oeb[PIN_VGA_VSYNC] = 1'b0;
	
	// IO37-PIN_VGA_HSYNC: Output
	localparam PIN_VGA_HSYNC = 37;
	assign gpio_input[PIN_VGA_HSYNC] = 1'b0;
	assign io_out[PIN_VGA_HSYNC] = vga_hsync;
	assign io_oeb[PIN_VGA_HSYNC] = 1'b0;
	
	//--------------End of Generated Code--------------//
	//-----------------Pin Mapping End-----------------//
	//-------------------------------------------------//

endmodulemodule PWM #(
		parameter ID = 8'h02
	)(

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		input wire clk,
		input wire rst,
		
		// Peripheral Bus
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[23:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,

		output wire[15:0] pwm_en,
		output wire[15:0] pwm_out,
		output wire[3:0] pwm_irq
	);

	localparam DEVICE_COUNT = 4;
	localparam OUTPUTS_PER_DEVICE = 4;

	// Peripheral select
	wire[15:0] localAddress;
	wire peripheralEnable;
	PeripheralSelect #(.ID(ID)) select(
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.peripheralEnable(peripheralEnable));
	
	wire[DEVICE_COUNT-1:0] deviceOutputRequest;
	wire[(32 * DEVICE_COUNT) - 1:0] deviceOutputData;
	Mux #(.WIDTH(32), .INPUTS(DEVICE_COUNT), .DEFAULT(~32'b0)) mux(
		.select(deviceOutputRequest),
		.in(deviceOutputData),
		.out(peripheralBus_dataRead),
		.outputEnable(requestOutput));

	wire[DEVICE_COUNT-1:0] deviceBusy_nc;

	genvar i;
	generate
		for (i = 0; i < DEVICE_COUNT; i = i + 1) begin			
			PWMDevice #(.ID(i+1), .OUTPUTS(OUTPUTS_PER_DEVICE), .WIDTH(16), .CLOCK_WIDTH(32)) device(
				.clk(clk),
				.rst(rst),
				.peripheralEnable(peripheralEnable),
				.peripheralBus_we(peripheralBus_we),
				.peripheralBus_oe(peripheralBus_oe),
				.peripheralBus_busy(deviceBusy_nc[i]),
				.peripheralBus_address(localAddress),
				.peripheralBus_byteSelect(peripheralBus_byteSelect),
				.peripheralBus_dataWrite(peripheralBus_dataWrite),
				.peripheralBus_dataRead(deviceOutputData[(i * 32) + 31:i * 32]),
				.requestOutput(deviceOutputRequest[i]),
				.pwm_en(pwm_en[(i * OUTPUTS_PER_DEVICE) + OUTPUTS_PER_DEVICE - 1:i * OUTPUTS_PER_DEVICE]),
				.pwm_out(pwm_out[(i * OUTPUTS_PER_DEVICE) + OUTPUTS_PER_DEVICE - 1:i * OUTPUTS_PER_DEVICE]),
				.pwm_irq(pwm_irq[i]));
		end
	endgenerate

	assign peripheralBus_busy = 1'b0;

endmodulemodule PWMDevice #(
		parameter ID = 4'h0,
		parameter OUTPUTS = 4,
		parameter WIDTH = 16,
		parameter CLOCK_WIDTH = 32
	)(
		input wire clk,
		input wire rst,

		// Peripheral bus
		input wire peripheralEnable,
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[15:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output reg[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,
		
		// PWM output
		output wire[OUTPUTS-1:0] pwm_en,
		output wire[OUTPUTS-1:0] pwm_out,
		output wire pwm_irq
	);

	localparam CLOCK_BITS = $clog2(CLOCK_WIDTH);

	wire counterEnable;
	wire[CLOCK_BITS-1:0] clockScale;
	wire[OUTPUTS-1:0] compareEnable;
	wire[OUTPUTS-1:0] outputEnable;
	wire[OUTPUTS-1:0] riseInterruptEnable;
	wire[OUTPUTS-1:0] fallInterruptEnable;

	// Counter control
	reg[CLOCK_WIDTH + WIDTH - 1:0] baseCounter = 'b0;
	wire[CLOCK_WIDTH + WIDTH - 1:0] nextCounter = baseCounter + 1;
	wire[WIDTH-1:0] counterValue = baseCounter >> clockScale;

	// Device select
	wire[11:0] localAddress;
	wire deviceEnable;
	DeviceSelect #(.ID(ID)) select(
		.peripheralEnable(peripheralEnable),
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.deviceEnable(deviceEnable));

	// Register
	// Configuration register 	 Default 0x000003 (for .CLOCK_WIDTH(32))
	// b00-b04: clockScale		 Default 0x03
	// b05: counterEnable		 Default 0x0
	// b06: compareEnable0		 Default 0x0
	// b07: compareEnable1		 Default 0x0
	// b08: compareEnable2		 Default 0x0
	// b09: compareEnable3		 Default 0x0
	// b10: outputEnable0		 Default 0x0
	// b11: outputEnable1		 Default 0x0
	// b12: outputEnable2		 Default 0x0
	// b13: outputEnable3		 Default 0x0
	// b14: riseInterruptEnable0 Default 0x0
	// b15: riseInterruptEnable1 Default 0x0
	// b16: riseInterruptEnable2 Default 0x0
	// b17: riseInterruptEnable3 Default 0x0
	// b18: fallInterruptEnable0 Default 0x0
	// b19: fallInterruptEnable1 Default 0x0
	// b20: fallInterruptEnable2 Default 0x0
	// b21: fallInterruptEnable3 Default 0x0
	localparam CONFIG_WIDTH = 1 + CLOCK_BITS + (OUTPUTS * 4);
	wire[CONFIG_WIDTH-1:0] configuration;
	wire[31:0] configurationRegisterOutputData;
	wire configurationRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(CONFIG_WIDTH), .ADDRESS(12'h000), .DEFAULT({ {(CONFIG_WIDTH-5){1'b0}}, 5'h0E })) configurationRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(configurationRegisterOutputData),
		.requestOutput(configurationRegisterOutputRequest),
		.currentValue(configuration));

	assign clockScale = configuration[CLOCK_BITS-1:0];
	assign counterEnable = configuration[CLOCK_BITS];
	assign compareEnable = configuration[(1 + CLOCK_BITS + OUTPUTS)-1:1 + CLOCK_BITS];
	assign outputEnable = configuration[(1 + CLOCK_BITS + (OUTPUTS * 2))-1:1 + CLOCK_BITS + OUTPUTS];
	assign riseInterruptEnable = configuration[(1 + CLOCK_BITS + (OUTPUTS * 3))-1:1 + CLOCK_BITS + (OUTPUTS * 2)];
	assign fallInterruptEnable = configuration[(1 + CLOCK_BITS + (OUTPUTS * 4))-1:1 + CLOCK_BITS + (OUTPUTS * 3)];

	// Counter top compare Default 0x1387 (for .WIDTH(16))
	// With clockScale=0x03, this gives a 1kHz signal with a 200ns resolution
	localparam DEFAULT_TOP_COMPARE_VALUE = 'h1387;
	wire[31:0] topCompareRegisterOutputData;
	wire topCompareRegisterOutputRequest;
	wire topCompareRegisterBusBusy_nc;
	wire[WIDTH-1:0] topCompareRegisterWriteData;
	wire topCompareRegisterWriteDataEnable;
	wire topCompareRegisterReadDataEnable_nc;
	reg[WIDTH-1:0] topCompare;
	DataRegister #(.WIDTH(WIDTH), .ADDRESS(12'h004)) topCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(topCompareRegisterBusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(topCompareRegisterOutputData),
		.requestOutput(topCompareRegisterOutputRequest),
		.writeData(topCompareRegisterWriteData),
		.writeData_en(topCompareRegisterWriteDataEnable),
		.writeData_busy(1'b0),
		.readData(topCompare),
		.readData_en(topCompareRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	// Current data register (for .WIDTH(16), .OUTPUTS(4))
	// b00-b15: counterValue
	// b16-b19: output
	reg[WIDTH+OUTPUTS-1:0] dataRegisterBuffered;
	wire[OUTPUTS-1:0] outputs;
	wire[31:0] dataRegisterOutputData;
	wire dataRegisterOutputRequest;
	wire dataRegisterBusBusy_nc;
	wire[WIDTH+OUTPUTS-1:0] dataRegisterWriteData_nc;
	wire dataRegisterWriteDataEnable_nc;
	wire dataRegisterReadDataEnable_nc;
	DataRegister #(.WIDTH(WIDTH + OUTPUTS), .ADDRESS(12'h008)) dataRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(dataRegisterBusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(dataRegisterOutputData),
		.requestOutput(dataRegisterOutputRequest),
		.writeData(dataRegisterWriteData_nc),
		.writeData_en(dataRegisterWriteDataEnable_nc),
		.writeData_busy(1'b0),
		.readData(dataRegisterBuffered),
		.readData_en(dataRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	always @(posedge clk) begin
		if (rst) dataRegisterBuffered <= {(WIDTH + OUTPUTS){1'b0}};
		else dataRegisterBuffered <= { outputs, counterValue };
	end

	always @(posedge clk) begin
		if (rst) begin
			baseCounter <= 'b0;
			topCompare <= DEFAULT_TOP_COMPARE_VALUE;
		end else begin
			if (topCompareRegisterWriteDataEnable) begin
				baseCounter <= 'b0;
				topCompare <= topCompareRegisterWriteData;
			end else begin
				if (counterEnable) begin
					if (counterValue == topCompare) baseCounter <= 'b0;
					else baseCounter <= nextCounter;
				end else begin
					baseCounter <= 'b0;
				end
			end
		end
	end

	wire[OUTPUTS-1:0] compareRegisterOutputRequest;
	wire[(32 * OUTPUTS) - 1:0] compareRegisterOutputData;
	wire[31:0] compareValuesOutputData;
	wire compareValuesOutputRequest;
	Mux #(.WIDTH(32), .INPUTS(OUTPUTS), .DEFAULT(~32'b0)) mux(
		.select(compareRegisterOutputRequest),
		.in(compareRegisterOutputData),
		.out(compareValuesOutputData),
		.outputEnable(compareValuesOutputRequest));

	assign requestOutput = configurationRegisterOutputRequest || topCompareRegisterOutputRequest || dataRegisterOutputRequest || compareValuesOutputRequest;

	always @(*) begin
		case (1'b1)
			configurationRegisterOutputRequest: peripheralBus_dataRead <= configurationRegisterOutputData;
			topCompareRegisterOutputRequest: peripheralBus_dataRead <= topCompareRegisterOutputData;
			dataRegisterOutputRequest: peripheralBus_dataRead <= dataRegisterOutputData;
			compareValuesOutputRequest: peripheralBus_dataRead <= compareValuesOutputData;
			default: peripheralBus_dataRead <= 32'b0;
		endcase
	end

	wire[OUTPUTS-1:0] compareRise;
	wire[OUTPUTS-1:0] compareFall;

	// Outputs
	genvar i;
	generate
		for (i = 0; i < OUTPUTS; i = i + 1) begin
			// Compare value register
			wire[WIDTH-1:0] compareValue;
			ConfigurationRegister #(.WIDTH(WIDTH), .ADDRESS(12'h010 + (i * 12'h004)), .DEFAULT('b0)) compareRegister(
				.clk(clk),
				.rst(rst),
				.enable(deviceEnable),
				.peripheralBus_we(peripheralBus_we),
				.peripheralBus_oe(peripheralBus_oe),
				.peripheralBus_address(localAddress),
				.peripheralBus_byteSelect(peripheralBus_byteSelect),
				.peripheralBus_dataWrite(peripheralBus_dataWrite),
				.peripheralBus_dataRead(compareRegisterOutputData[(i * 32) + 31:i * 32]),
				.requestOutput(compareRegisterOutputRequest[i]),
				.currentValue(compareValue));
			PWMOutput #(.WIDTH(WIDTH)) outputPort(
				.clk(clk),
				.rst(rst),
				.compareValue(compareValue),
				.enable(compareEnable[i]),
				.counterValue(counterValue),
				.pwm_out(outputs[i]),
				.compareRise(compareRise[i]),
				.compareFall(compareFall[i]));
		end
	endgenerate

	assign peripheralBus_busy = 1'b0;

	assign pwm_en = compareEnable & outputEnable;
	assign pwm_out = outputs;

	wire[OUTPUTS-1:0] comparatorIRQ = (riseInterruptEnable & compareRise) || (fallInterruptEnable & compareFall);
	assign pwm_irq = |comparatorIRQ;

endmodule
module PWMOutput #(
		parameter WIDTH = 16
	)(
		input wire clk,
		input wire rst,
		
		input wire[WIDTH-1:0] compareValue,
		input wire enable,

		input wire[WIDTH-1:0] counterValue,
		output wire pwm_out,
		
		output reg compareRise,
		output reg compareFall
	);

	reg [WIDTH-1:0] currentCompareValue = {WIDTH{1'b0}};
	wire equality = counterValue == currentCompareValue;

	reg state = 1'b0;

	always @(posedge clk) begin
		if (rst) begin
			currentCompareValue <= {WIDTH{1'b0}};
			state <= 1'b0;
		end else begin
			if (enable) begin
				if (counterValue == 0) begin
					state <= 1'b0;
					currentCompareValue <= compareValue;
				end	else if (equality) begin
					state <= 1'b1;
				end
			end else begin
				state <= 1'b0;
				currentCompareValue <= compareValue;
			end
		end
	end

	reg lastState = 1'b0;
	always @(posedge clk) begin
		if (rst) begin
			lastState <= 1'b0;
			compareRise <= 1'b0;
			compareFall <= 1'b0;
		end	else begin 
			lastState <= state;

			if (state != state) begin
				compareRise <= state;
				compareFall <= !state;
			end else begin
				compareRise <= 1'b0;
				compareFall <= 1'b0;
			end
		end
	end
	
	assign pwm_out = state;

endmodulemodule SPI #(
		parameter ID = 8'h01
	)(

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		input wire clk,
		input wire rst,
		
		// Peripheral Bus
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[23:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,

		output wire[DEVICE_COUNT-1:0] spi_en,
		output wire[DEVICE_COUNT-1:0] spi_clk,
		output wire[DEVICE_COUNT-1:0] spi_mosi,
		input  wire[DEVICE_COUNT-1:0] spi_miso,
		output wire[DEVICE_COUNT-1:0] spi_cs
	);

	localparam DEVICE_COUNT = 1;

	// Peripheral select
	wire[15:0] localAddress;
	wire peripheralEnable;
	PeripheralSelect #(.ID(ID)) select(
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.peripheralEnable(peripheralEnable));

	wire[DEVICE_COUNT-1:0] deviceBusy;
	wire[DEVICE_COUNT-1:0] deviceOutputRequest;
	wire[(32 * DEVICE_COUNT) - 1:0] deviceOutputData;
	Mux #(.WIDTH(32), .INPUTS(DEVICE_COUNT), .DEFAULT(~32'b0)) mux(
		.select(deviceOutputRequest),
		.in(deviceOutputData),
		.out(peripheralBus_dataRead),
		.outputEnable(requestOutput));

	genvar i;
	generate
		for (i = 0; i < DEVICE_COUNT; i = i + 1) begin
			SPIDevice #(.ID(i+1), .CLOCK_WIDTH(8)) device(
				.clk(clk),
				.rst(rst),
				.peripheralEnable(peripheralEnable),
				.peripheralBus_we(peripheralBus_we),
				.peripheralBus_oe(peripheralBus_oe),
				.peripheralBus_busy(deviceBusy[i]),
				.peripheralBus_address(localAddress),
				.peripheralBus_byteSelect(peripheralBus_byteSelect),
				.peripheralBus_dataWrite(peripheralBus_dataWrite),
				.peripheralBus_dataRead(deviceOutputData[(i * 32) + 31:i * 32]),
				.requestOutput(deviceOutputRequest[i]),
				.spi_en(spi_en[i]),
				.spi_clk(spi_clk[i]),
				.spi_mosi(spi_mosi[i]),
				.spi_miso(spi_miso[i]),
				.spi_cs(spi_cs[i]));
		end
	endgenerate
	
	assign peripheralBus_busy = |deviceBusy;

endmodulemodule SPIDevice #(
		parameter ID = 4'h0,
		parameter CLOCK_WIDTH = 8
	)(
		input wire clk,
		input wire rst,

		// Peripheral bus
		input wire peripheralEnable,
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[15:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output reg[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,

		// SPI interface
		output wire spi_en,
		output reg spi_clk,
		output wire spi_mosi,
		input  wire spi_miso,
		output wire spi_cs
	);

	localparam CLOCK_BITS = $clog2(CLOCK_WIDTH);

	localparam STATE_IDLE  = 2'b00;
	localparam STATE_SETUP = 2'b01;
	localparam STATE_SHIFT = 2'b10;
	localparam STATE_END   = 2'b11;

	// Device select
	wire[11:0] localAddress;
	wire deviceEnable;
	DeviceSelect #(.ID(ID)) select(
		.peripheralEnable(peripheralEnable),
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.deviceEnable(deviceEnable));

	// Register
	// Configuration register 	Default 0x064
	// b00-b02: clockScale 		Default 0x4
	// b03-04: spiMode 			Default 0x0
	// b05: msbFirst 			Default 0x1
	// b06: useCS 				Default 0x1
	// b07: activeHighCS		Default 0x0
	// b08: enable				Default 0x0
	wire[31:0] configurationRegisterOutputData;
	wire configurationRegisterOutputRequest;
	wire[8:0] configuration;
	ConfigurationRegister #(.WIDTH(9), .ADDRESS(12'h000), .DEFAULT(9'h064)) configurationRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(configurationRegisterOutputData),
		.requestOutput(configurationRegisterOutputRequest),
		.currentValue(configuration));

	wire[2:0] clockScale = configuration[2:0];
	wire[1:0] spiMode = configuration[4:3];
	wire msbFirst = configuration[5];
	wire useCS = configuration[6];
	wire activeHighCS = configuration[7];
	assign spi_en = configuration[8];
	wire spiClockPolarity = spiMode[1];
	wire spiSampleMode = spiMode[0];

	// Status register
	wire deviceBusy = state != STATE_IDLE;
	wire[31:0] statusRegisterOutputData;
	wire statusRegisterOutputRequest;
	wire statusRegisterWriteData_nc;
	wire statusRegisterWriteDataEnable_nc;
	wire statusRegisterReadDataEnable_nc;
	wire statusRegisterBusBusy_nc;
	DataRegister #(.WIDTH(1), .ADDRESS(12'h004)) statusRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(statusRegisterBusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(statusRegisterOutputData),
		.requestOutput(statusRegisterOutputRequest),
		.writeData(statusRegisterWriteData_nc),
		.writeData_en(statusRegisterWriteDataEnable_nc),
		.writeData_busy(1'b0),
		.readData(deviceBusy),
		.readData_en(statusRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	// Input and Output register
	wire[31:0] dataRegisterOutputData;
	wire dataRegisterOutputRequest;
	wire[7:0] dataRegisterReadData;
	wire[7:0] dataRegisterWriteData;	
	wire dataRegisterWriteDataEnable;
	wire dataRegisterBusBusy;
	wire dataRegisterReadDataEnable_nc;
	DataRegister #(.WIDTH(8), .ADDRESS(12'h008)) dataRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(dataRegisterBusBusy),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(dataRegisterOutputData),
		.requestOutput(dataRegisterOutputRequest),
		.writeData(dataRegisterWriteData),
		.writeData_en(dataRegisterWriteDataEnable),
		.writeData_busy(deviceBusy),
		.readData(dataRegisterReadData),
		.readData_en(dataRegisterReadDataEnable_nc),
		.readData_busy(deviceBusy));

	// State control
	reg[1:0] state = STATE_IDLE;
	
	reg[2:0] bitCounter = 3'b0;
	wire[2:0] nextBitCounter = bitCounter + 1;

	reg[CLOCK_WIDTH-1:0] clockCounter = {CLOCK_WIDTH{1'b0}};
	wire[CLOCK_WIDTH-1:0] nextClockCounter = clockCounter + 1;
	wire[CLOCK_WIDTH-1:0] clockScaleCompare = { {(CLOCK_WIDTH-1){1'b0}}, 1'b1 } << clockScale;
	wire[CLOCK_WIDTH-1:0] clockScaleHalfCompare = { 1'b0, clockScaleCompare[CLOCK_WIDTH-1:1] };
	wire halfClockCounterMatch = nextClockCounter == clockScaleHalfCompare;
	wire clockCounterMatch     = nextClockCounter == clockScaleCompare;

	reg spiClockRise = 1'b0;
	reg spiClockFall = 1'b0;
	reg spiClock;

	wire shiftInEnable  = spiSampleMode ? spiClockFall : spiClockRise;
	wire shiftOutEnable = spiSampleMode ? spiClockRise : spiClockFall;
	
	wire serialOut;
	ShiftRegister #(.WIDTH(8)) register (
		.clk(clk),
		.rst(rst),
		.loadEnable(dataRegisterWriteDataEnable),
		.shiftInEnable(shiftInEnable),
		.shiftOutEnable(shiftOutEnable),
		.msbFirst(msbFirst),
		.parallelIn(dataRegisterWriteData),
		.parallelOut(dataRegisterReadData),
		.serialIn(spi_miso),
		.serialOut(serialOut));

	always @(posedge clk) begin
		if (rst) begin
			state <= STATE_IDLE;
			bitCounter <= 3'b0;
			clockCounter <= {CLOCK_WIDTH{1'b0}};
			spiClockRise <= 1'b0;
			spiClockFall <= 1'b0;
			spiClock <= 1'b0;
		end else begin
			case (state)
				STATE_IDLE: begin
					bitCounter <= 3'b0;
					clockCounter <= {CLOCK_WIDTH{1'b0}};
					spiClockRise <= 1'b0;
					spiClockFall <= 1'b0;
					spiClock <= 1'b0;

					if (dataRegisterWriteDataEnable && peripheralBus_byteSelect[0]) begin 
						state <= STATE_SETUP;
					end
				end

				STATE_SETUP: begin
					clockCounter <= nextClockCounter;

					if (halfClockCounterMatch) begin
						bitCounter <= 1'b0;
						spiClock <= 1'b1;
						state <= STATE_SHIFT;

						if (spiClockPolarity) begin
							spiClockRise <= 1'b0;
							spiClockFall <= 1'b1;
						end else begin
							spiClockRise <= 1'b1;
							spiClockFall <= 1'b0;
						end	
					end					
				end

				STATE_SHIFT: begin
					if (clockCounterMatch) begin
						clockCounter <= {CLOCK_WIDTH{1'b0}};
						spiClock <= 1'b0;

						if (spiClockPolarity) begin
							spiClockRise <= 1'b1;
							spiClockFall <= 1'b0;
						end else begin
							spiClockRise <= 1'b0;
							spiClockFall <= 1'b1;
						end

						if (bitCounter == 3'h7) begin
							state <= STATE_END;
						end	else begin
							bitCounter <= nextBitCounter;
						end
					end else if (halfClockCounterMatch) begin
						if (spiClockPolarity) begin
							spiClockRise <= 1'b0;
							spiClockFall <= 1'b1;
						end else begin
							spiClockRise <= 1'b1;
							spiClockFall <= 1'b0;
						end	

						spiClock <= 1'b1;
						clockCounter <= nextClockCounter;
					end else begin
						spiClockRise <= 1'b0;
						spiClockFall <= 1'b0;
						clockCounter <= nextClockCounter;
					end
				end

				STATE_END: begin
					spiClockRise <= 1'b0;
					spiClockFall <= 1'b0;
					spiClock <= 1'b0;
					
					if (clockCounterMatch) state <= STATE_IDLE;
					else clockCounter <= nextClockCounter;
				end

				default: begin
					state <= STATE_IDLE;
					bitCounter <= 3'b0;
					clockCounter <= {CLOCK_WIDTH{1'b0}};
					spiClockRise <= 1'b0;
					spiClockFall <= 1'b0;
					spiClock <= 1'b0;
				end
			endcase
		end
	end

	// Buffer the spi clock by one cycle so that it lines up with when data is sampled
	always @(posedge clk) begin
		if (rst) spi_clk <= 1'b0;
		else spi_clk <= spiClockPolarity ? !spiClock : spiClock;
	end

	assign requestOutput = configurationRegisterOutputRequest || statusRegisterOutputRequest || dataRegisterOutputRequest;

	always @(*) begin
		case (1'b1)
			configurationRegisterOutputRequest: peripheralBus_dataRead <= configurationRegisterOutputData;
			statusRegisterOutputRequest: peripheralBus_dataRead <= statusRegisterOutputData;
			dataRegisterOutputRequest: peripheralBus_dataRead <= dataRegisterOutputData;
			default: peripheralBus_dataRead <=  ~32'b0;
		endcase
	end

	assign peripheralBus_busy = dataRegisterBusBusy;

	assign spi_mosi = serialOut & deviceBusy;
	assign spi_cs = useCS ? (activeHighCS ? deviceBusy : !deviceBusy) : 1'b0;

endmodulemodule UART #(
		parameter ID = 8'h00
	)(

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		input wire clk,
		input wire rst,
		
		// Peripheral Bus
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[23:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,

		// UART
		output wire[3:0] uart_en,	
		input wire[3:0] uart_rx,
		output wire[3:0] uart_tx,
		output wire[3:0] uart_irq
	);

	localparam DEVICE_COUNT = 4;

	// Peripheral select
	wire[15:0] localAddress;
	wire peripheralEnable;
	PeripheralSelect #(.ID(ID)) select(
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.peripheralEnable(peripheralEnable));

	wire[DEVICE_COUNT-1:0] deviceBusy;
	wire[DEVICE_COUNT-1:0] deviceOutputRequest;
	wire[(32 * DEVICE_COUNT) - 1:0] deviceOutputData;
	Mux #(.WIDTH(32), .INPUTS(DEVICE_COUNT), .DEFAULT(~32'b0)) mux(
		.select(deviceOutputRequest),
		.in(deviceOutputData),
		.out(peripheralBus_dataRead),
		.outputEnable(requestOutput));

	genvar i;
	generate
		for (i = 0; i < DEVICE_COUNT; i = i + 1) begin
			UARTDevice #(.ID(i+1)) device(
				.clk(clk),
				.rst(rst),
				.peripheralEnable(peripheralEnable),
				.peripheralBus_we(peripheralBus_we),
				.peripheralBus_oe(peripheralBus_oe),
				.peripheralBus_busy(deviceBusy[i]),
				.peripheralBus_address(localAddress),
				.peripheralBus_byteSelect(peripheralBus_byteSelect),
				.peripheralBus_dataWrite(peripheralBus_dataWrite),
				.peripheralBus_dataRead(deviceOutputData[(i * 32) + 31:i * 32]),
				.requestOutput(deviceOutputRequest[i]),
				.uart_en(uart_en[i]),
				.uart_rx(uart_rx[i]),
				.uart_tx(uart_tx[i]),
				.uart_irq(uart_irq[i]));
		end
	endgenerate

	assign peripheralBus_busy = |deviceBusy;

endmodulemodule UARTDevice  #(
		parameter ID = 4'h0
	)(
		input wire clk,
		input wire rst,

		// Peripheral bus
		input wire peripheralEnable,
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[15:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,
		
		// PWM output
		output wire uart_en,
		input wire uart_rx,
		output wire uart_tx,
		output wire uart_irq
	);

	localparam RX_BUFFER_SIZE = 32;
	localparam TX_BUFFER_SIZE = 32;

	// Buffer values used for interrupts and status register
	wire txDataLost;
	wire txBufferFull;
	wire txDataAvailable;
	wire rxDataLost;
	wire rxBufferFull;
	wire rxDataAvailable;

	reg txDataLostBuffered;
	reg txBufferFullBuffered;
	reg txDataAvailableBuffered;
	reg rxDataLostBuffered;
	reg rxBufferFullBuffered;
	reg rxDataAvailableBuffered;

	always @(posedge clk) begin
		if (rst) begin
			txDataLostBuffered <= 1'b0;
			txBufferFullBuffered <= 1'b0;
			txDataAvailableBuffered <= 1'b0;
			rxDataLostBuffered <= 1'b0;
			rxBufferFullBuffered <= 1'b0;
			rxDataAvailableBuffered <= 1'b0;
		end else begin
			txDataLostBuffered <= txDataLost;
			txBufferFullBuffered <= txBufferFull;
			txDataAvailableBuffered <= txDataAvailable;
			rxDataLostBuffered <= rxDataLost;
			rxBufferFullBuffered <= rxBufferFull;
			rxDataAvailableBuffered <= rxDataAvailable;
		end
	end

	// Device select
	wire[11:0] localAddress;
	wire deviceEnable;
	DeviceSelect #(.ID(ID)) select(
		.peripheralEnable(peripheralEnable),
		.peripheralBus_address(peripheralBus_address),
		.localAddress(localAddress),
		.deviceEnable(deviceEnable));

	// Register
	// Configuration register 				Default 0x01047
	// b00-b15: cyclesPerBit  				Default 0x1047	((CLK_FREQ + BAUD) / BAUD) - 1 => Default uses CLK_FREQ=40MHz BAUD=9600(Actually 9599.2)
	// b16: waitForTxSpace	  				Default 0x0
	// b17: enable 			  				Default 0x0
	// b18: dataLostInterruptEnable			Default 0x0
	// b19: rxDataAvaliableInterruptEnable	Default 0x0
	// b20: txDataSentInterruptEnable		Default 0x0
	wire[31:0] configurationRegisterOutputData;
	wire configurationRegisterOutputRequest;
	wire[20:0] configuration;
	ConfigurationRegister #(.WIDTH(21), .ADDRESS(12'h000), .DEFAULT(21'h001047)) configurationRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(configurationRegisterOutputData),
		.requestOutput(configurationRegisterOutputRequest),
		.currentValue(configuration));

	wire[15:0] cyclesPerBit = configuration[15:0];
	wire waitForTxSpace = configuration[16];
	assign uart_en = configuration[17];
	wire dataLostInterruptEnable = configuration[18];
	wire rxDataAvaliableInterruptEnable = configuration[19];
	wire txDataSentInterruptEnable = configuration[20];

	// Clear register
	wire[3:0] clearWriteData;
	wire clearWriteEnable;
	wire clearRegisterBusyBusy_nc;
	wire[31:0] clearRegisterDataOut;
	wire clearRegisterRequestOutput_nc;
	wire clearRegisterReadDataEnable_nc;
	DataRegister #(.WIDTH(4), .ADDRESS(12'h004)) clearRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(clearRegisterBusyBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(clearRegisterDataOut),
		.requestOutput(clearRegisterRequestOutput_nc),
		.writeData(clearWriteData),
		.writeData_en(clearWriteEnable),
		.writeData_busy(1'b0),
		.readData(4'b0),
		.readData_en(clearRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	// Status register
	// b00: rxDataAvailable
	// b01: rxBufferFull
	// b02: rxDataLost
	// b03: txDataAvailable
	// b04: txBufferFull
	// b05: txDataLost
	reg[5:0] statusRegisterBuffered;
	wire[31:0] statusRegisterOutputData;
	wire statusRegisterOutputRequest;
	wire statusRegisterBusBusy_nc;
	wire[5:0] statusRegisterWriteData_nc;
	wire statusRegisterWriteDataEnable_nc;
	wire statusRegisterReadDataEnable_nc;
	DataRegister #(.WIDTH(6), .ADDRESS(12'h008)) statusRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(statusRegisterBusBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(statusRegisterOutputData),
		.requestOutput(statusRegisterOutputRequest),
		.writeData(statusRegisterWriteData_nc),
		.writeData_en(statusRegisterWriteDataEnable_nc),
		.writeData_busy(1'b0),
		.readData(statusRegisterBuffered),
		.readData_en(statusRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	always @(posedge clk) begin
		if (rst) statusRegisterBuffered <= 6'b0;
		else begin
			statusRegisterBuffered <= { 
				txDataLostBuffered, 
				txBufferFullBuffered, 
				txDataAvailableBuffered, 
				rxDataLostBuffered, 
				rxBufferFullBuffered, 
				rxDataAvailableBuffered
			};
		end
	end

	// Rx register
	reg[8:0] rxRegisterBuffered;
	wire[31:0] rxRegisterOutputData;
	wire rxRegisterOutputRequest;
	wire[7:0] rxReadData;
	wire rxReadDataEnable;
	wire rxRegisterBusyBusy_nc;
	wire[8:0] rxRegisterWriteData_nc;
	wire rxRegisterWriteDataEnable_nc;
	DataRegister #(.WIDTH(9), .ADDRESS(12'h010)) rxRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(rxRegisterBusyBusy_nc),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(rxRegisterOutputData),
		.requestOutput(rxRegisterOutputRequest),
		.writeData(rxRegisterWriteData_nc),
		.writeData_en(rxRegisterWriteDataEnable_nc),
		.writeData_busy(1'b0),
		.readData(rxRegisterBuffered),
		.readData_en(rxReadDataEnable),
		.readData_busy(1'b0));

	always @(posedge clk) begin
		if (rst) rxRegisterBuffered <= 9'b0;
		else rxRegisterBuffered <= rxDataAvailable ? { 1'b1, rxReadData } : 9'h0;
	end

	// Tx register
	wire[31:0] txRegisterOutputData;
	wire txRegisterOutputRequest;
	wire[7:0] txWriteData;	
	wire txWriteDataEnable;
	wire txBusy;
	wire txRegisterReadDataEnable_nc;
	DataRegister #(.WIDTH(8), .ADDRESS(12'h014)) txRegister(
		.clk(clk),
		.rst(rst),
		.enable(deviceEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(txBusy),
		.peripheralBus_address(localAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(txRegisterOutputData),
		.requestOutput(txRegisterOutputRequest),
		.writeData(txWriteData),
		.writeData_en(txWriteDataEnable),
		.writeData_busy(waitForTxSpace && txBufferFull && uart_en),
		.readData(8'b0),
		.readData_en(txRegisterReadDataEnable_nc),
		.readData_busy(1'b0));

	wire [7:0] rxByteIn;
	wire rxOutAvailable;
	UART_rx #(.CLOCK_SCALE_BITS(16)) uartRx(
		.clk(clk),
		.rst(rst || (clearWriteData[0] && clearWriteEnable && peripheralBus_byteSelect[0])),
		.cyclesPerBit(cyclesPerBit),
		.rx(uart_en ? uart_rx : 1'b1),
		.dataOut(rxByteIn),
		.dataAvailable(rxOutAvailable));
	
	wire txSendBusy;
	wire[7:0] txByteOut;
	UART_tx #(.CLOCK_SCALE_BITS(16)) uartTx(
		.clk(clk),
		.rst(rst || (clearWriteData[1] && clearWriteEnable && peripheralBus_byteSelect[0])),
		.cyclesPerBit(cyclesPerBit),
		.tx(uart_tx),
		.blockTransmition(!uart_en),
    	.busy(txSendBusy),
    	.dataIn(txByteOut),
    	.dataAvailable(txDataAvailable));

	FIFO #(.WORD_SIZE(8), .BUFFER_SIZE(RX_BUFFER_SIZE)) rxBuffer(
		.clk(clk),
		.rst(rst || (clearWriteData[2] && clearWriteEnable && peripheralBus_byteSelect[0])),
		.dataIn(rxByteIn),
		.we(rxOutAvailable && uart_en),
		.dataOut(rxReadData),
		.oe(rxReadDataEnable),		
		.isData(rxDataAvailable),
		.bufferFull(rxBufferFull),
		.dataLost(rxDataLost));

	FIFO #(.WORD_SIZE(8), .BUFFER_SIZE(TX_BUFFER_SIZE)) txBuffer(
		.clk(clk),
		.rst(rst || (clearWriteData[3] && clearWriteEnable && peripheralBus_byteSelect[0])),
		.dataIn(txWriteData),
		.we(txWriteDataEnable && peripheralBus_byteSelect[0] && (!waitForTxSpace || !txBufferFull)),
		.dataOut(txByteOut),
		.oe(txDataAvailable && uart_en && !txSendBusy),		
		.isData(txDataAvailable),
		.bufferFull(txBufferFull),
		.dataLost(txDataLost));

	assign requestOutput = configurationRegisterOutputRequest || statusRegisterOutputRequest || rxRegisterOutputRequest || txRegisterOutputRequest;
	assign peripheralBus_dataRead = configurationRegisterOutputRequest ? configurationRegisterOutputData :
									statusRegisterOutputRequest		   ? statusRegisterOutputData :
								    rxRegisterOutputRequest 		   ? rxRegisterOutputData :
									txRegisterOutputRequest 		   ? txRegisterOutputData :
													   					 ~32'b0;
	assign peripheralBus_busy = txBusy;

	reg sendingData = 1'b0;
	always @(posedge clk) begin
		if (rst) sendingData <= 1'b0;
		else sendingData <= txDataAvailableBuffered;
	end

	assign uart_irq = (dataLostInterruptEnable && (rxDataLostBuffered || txDataLostBuffered))
				   || (rxDataAvaliableInterruptEnable && rxDataAvailableBuffered)
				   || (txDataSentInterruptEnable && sendingData && !txDataAvailableBuffered);

endmodulemodule UART_rx
	#(
		parameter CLOCK_SCALE_BITS = 16
	)(
		input wire clk,
		input wire rst,
		input wire[CLOCK_SCALE_BITS-1:0] cyclesPerBit, // ((CLK_FREQ + BAUD) / BAUD) - 1
		input wire rx,
		output wire [7:0] dataOut,
    	output wire dataAvailable
    );

	localparam STATE_IDLE		= 2'b00;
	localparam STATE_WAIT_HALF 	= 2'b01;
	localparam STATE_WAIT_FULL 	= 2'b10;
	localparam STATE_WAIT_HIGH 	= 2'b11;

	reg[1:0] state = STATE_IDLE;
	reg[CLOCK_SCALE_BITS-1:0] delayCounter = {CLOCK_SCALE_BITS{1'b0}};
	wire[CLOCK_SCALE_BITS-1:0] nextDelayCounter = delayCounter + 1;

	reg[2:0] bitCounter = 3'b0;
	reg[7:0] savedData = 8'b0;
	reg newData = 1'b0;

	wire[CLOCK_SCALE_BITS-1:0] halfBitCounterValue = { 1'b0, cyclesPerBit[CLOCK_SCALE_BITS-1:1] };

	always @(posedge clk) begin
		if (rst) begin
			state = STATE_IDLE;
			delayCounter = {CLOCK_SCALE_BITS{1'b0}};
			bitCounter = 3'b0;
			savedData = 8'b0;
			newData = 1'b0;
		end else begin
			newData = 1'b0;

			 /* When a new byte is being received, the input goes low. This is the
				start bit. When the beginning of this bit is detected we need to wait
				one and a half bit widths before reading in the first data bit. The
				half cycle is so that we read in the middle of the bit for the most
				accurate result. WAIT_HALF waits this half cycle and WAIT_FULL waits
				a full cycle then reads in a bit. After 8 bits are read, the data is
				output and the FSM waits for the RX input to go high again to signal
				the end of the transmission. The FSM then returns to IDLE ready to
				receive the next byte.                                               */
			case (state)
				STATE_IDLE: begin
					bitCounter = 3'b0;
					delayCounter = {CLOCK_SCALE_BITS{1'b0}};
					if (!rx) state = STATE_WAIT_HALF;
				end

				STATE_WAIT_HALF: begin
					if (nextDelayCounter == halfBitCounterValue) begin						
						delayCounter = 0;
						state = STATE_WAIT_FULL;
					end else begin
						delayCounter = nextDelayCounter;
					end
				end

				STATE_WAIT_FULL: begin
					if (nextDelayCounter == cyclesPerBit) begin
						savedData = {rx, savedData[7:1]};
						delayCounter = 0;
						if (bitCounter == 3'h7) begin
							state = STATE_WAIT_HIGH;
							newData = 1'b1;
						end else bitCounter = bitCounter + 1;
					end else begin
						delayCounter = nextDelayCounter;
					end
				end

				STATE_WAIT_HIGH: begin
					 if (rx) state = STATE_IDLE;
				end

				default: state = STATE_IDLE;				
			endcase
		end
	end

	assign dataOut = savedData;
	assign dataAvailable = newData;
endmodule
module UART_tx
	#(
		parameter CLOCK_SCALE_BITS = 16
	)(
		input wire clk,
		input wire rst,
		input wire[CLOCK_SCALE_BITS-1:0] cyclesPerBit, // ((CLK_FREQ + BAUD) / BAUD) - 1		
		output wire tx,
		input wire blockTransmition,
    	output reg busy,
    	input wire [7:0] dataIn,
    	input wire dataAvailable
    );
	
	localparam STATE_IDLE		= 2'b00;
	localparam STATE_START_BIT 	= 2'b01;
	localparam STATE_DATA 		= 2'b10;
	localparam STATE_STOP_BIT 	= 2'b11;

	reg[1:0] state = STATE_IDLE;
	reg[CLOCK_SCALE_BITS-1:0] delayCounter = {CLOCK_SCALE_BITS{1'b0}};
	wire[CLOCK_SCALE_BITS-1:0] nextDelayCounter = delayCounter + 1;
		
	reg[2:0] bitCounter = 3'b0;
	reg[7:0] savedData = 8'b0;
	reg outputBuffer = 1'b0;

	always @(posedge clk) begin
		if (rst) begin
			state = STATE_IDLE;
			delayCounter = {CLOCK_SCALE_BITS{1'b0}};
			bitCounter = 3'b0;
			savedData = 8'b0;
			outputBuffer = 1'b1;
		end else begin
			busy = 1'b1;
			
			/*  When a new byte is presnted to send, that byte is saved so that
				if the input changes the correct data is still sent. We first
				have to send a 0, which is the start bit. Once the start bit
				is sent, each data bit is sent out. The counter ctr is used to
				delay between bits to get the correct baud rate. The counter
				bitCounter is used to keep track of what bit to send. After
				all eight bits are sent, we need to send 1, the stop bit.
				This bit ensures that the line goes high between transmissions.
				When the transmistter is sending out data, the output busy is
				set to 1. To prevent the transmitter from sending data, set
				block to 1. This can be used for flow control.                  */
			case (state)
				STATE_IDLE: begin
					outputBuffer = 1'b1; // UART standard is to default to high

					if (!blockTransmition) begin
						busy = 1'b0;
						delayCounter = {CLOCK_SCALE_BITS{1'b0}};
						bitCounter = 3'b0;

						if (dataAvailable) begin
							savedData = dataIn;
							state = STATE_START_BIT;
						end
					end
				end

				STATE_START_BIT: begin
					outputBuffer = 1'b0;

					if (nextDelayCounter == cyclesPerBit) begin
						delayCounter = 0;
						state = STATE_DATA;
					end else begin
						delayCounter = nextDelayCounter;
					end
				end

				STATE_DATA: begin
					outputBuffer = savedData[bitCounter];

					if (nextDelayCounter == cyclesPerBit) begin
						delayCounter = 0;
						if (bitCounter == 3'h7) state = STATE_STOP_BIT;
						else bitCounter = bitCounter + 1;
					end else begin
						delayCounter = nextDelayCounter;
					end
				end

				STATE_STOP_BIT: begin
					outputBuffer = 1'b1;

					if (nextDelayCounter == cyclesPerBit) begin
						state = STATE_IDLE;
					end else begin
						delayCounter = nextDelayCounter;
					end
				end
				
				default: state = STATE_IDLE;				
			endcase
		end
	end

	assign tx = outputBuffer;

endmodule
module ConfigurationRegister #(
		parameter WIDTH = 32,
		parameter ADDRESS = 12'b0,
		parameter DEFAULT = 32'b0
	)(
		input wire clk,
		input wire rst,

		// Peripheral Bus
		input wire enable,
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		input wire[11:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,

		output wire[WIDTH-1:0] currentValue
	);
	
	wire[31:0] dataMask = {
		peripheralBus_byteSelect[3] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[2] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[1] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[0] ? 8'hFF : 8'h00
	};

	reg[WIDTH-1:0] registerValue;
	wire[31:0] maskedWriteData = (peripheralBus_dataWrite & dataMask) | (registerValue & ~dataMask);

	wire registerSelect = enable && ({ peripheralBus_address[11:2], 2'b00 } == ADDRESS);
	wire we = registerSelect && peripheralBus_we && !peripheralBus_oe;
	wire oe = registerSelect && peripheralBus_oe && !peripheralBus_we;

	always @(posedge clk) begin
		if (rst) begin
			registerValue <= DEFAULT;
		end else begin
			if (we) registerValue <= maskedWriteData[WIDTH-1:0];
		end
	end

	wire[31:0] baseReadData;
	generate
		if (WIDTH == 32) begin
			assign baseReadData = registerValue;
		end else begin
			wire[32-WIDTH-1:0] zeroPadding = 'b0;
			assign baseReadData = { zeroPadding, registerValue };
		end
	endgenerate

	assign peripheralBus_dataRead = oe ? baseReadData & dataMask : 32'b0;
	assign requestOutput = oe;
	assign currentValue = registerValue;

endmodulemodule DataRegister #(
		parameter WIDTH = 32,
		parameter ADDRESS = 12'b0
	)(
		input wire clk,
		input wire rst,

		// Peripheral Bus
		input wire enable,
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[11:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,

		output wire[WIDTH-1:0] writeData,
		output wire writeData_en,
		input wire writeData_busy,
		input wire[WIDTH-1:0] readData,
		output wire readData_en,
		input wire readData_busy
	);
	
	wire[31:0] dataMask = {
		peripheralBus_byteSelect[3] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[2] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[1] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[0] ? 8'hFF : 8'h00
	};

	wire registerSelect = enable && ({ peripheralBus_address[11:2], 2'b00 } == ADDRESS);
	wire we = registerSelect && peripheralBus_we && !peripheralBus_oe;
	wire oe = registerSelect && peripheralBus_oe && !peripheralBus_we;

	assign writeData = we ? peripheralBus_dataWrite[WIDTH-1:0] : {WIDTH{1'b0}};
	assign writeData_en = we;

	wire[31:0] baseReadData;
	generate
		if (WIDTH == 32) begin
			assign baseReadData = readData;
		end else begin
			wire[32-WIDTH-1:0] zeroPadding = 'b0;
			assign baseReadData = { zeroPadding, readData };
		end
	endgenerate

	assign peripheralBus_dataRead = oe ? baseReadData & dataMask : 32'b0;
	assign peripheralBus_busy = registerSelect && ((we && writeData_busy) | (oe && readData_busy));
	assign requestOutput = oe;
	assign readData_en = oe;

endmodulemodule OutputRegister #(
		parameter WIDTH = 32,
		parameter ADDRESS = 8'b0,
		parameter DEFAULT = 32'b0
	)(
		input wire clk,
		input wire rst,

		// Peripheral Bus
		input wire enable,
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		input wire[11:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		output wire[31:0] peripheralBus_dataRead,
		input wire[31:0] peripheralBus_dataWrite,
		output wire requestOutput,

		output wire[WIDTH-1:0] currentValue
	);
	
	localparam WRITE_ADDRESS = 4'h0;
	localparam SET_ADDRESS = 4'h4;
	localparam CLEAR_ADDRESS = 4'h8;
	localparam TOGGLE_ADDRESS = 4'hC;

	wire enableWrite = peripheralBus_address[3:0] == WRITE_ADDRESS;
	wire enableSet = peripheralBus_address[3:0] == SET_ADDRESS;
	wire enableClear = peripheralBus_address[3:0] == CLEAR_ADDRESS;
	wire enableToggle = peripheralBus_address[3:0] == TOGGLE_ADDRESS;

	wire[31:0] dataMask = {
		peripheralBus_byteSelect[3] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[2] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[1] ? 8'hFF : 8'h00,
		peripheralBus_byteSelect[0] ? 8'hFF : 8'h00
	};

	reg[WIDTH-1:0] registerValue;

	wire[31:0] maskedDataWrite = peripheralBus_dataWrite & dataMask;
	
	wire[31:0] writeData = maskedDataWrite | (registerValue & ~dataMask);
	wire[31:0] setData = registerValue | maskedDataWrite;
	wire[31:0] clearData = registerValue & ~maskedDataWrite;
	wire[31:0] toggleData = registerValue ^ maskedDataWrite;

	wire registerSelect = enable && (peripheralBus_address[11:4] == ADDRESS);
	wire we = registerSelect && peripheralBus_we && !peripheralBus_oe;
	wire oe = registerSelect && peripheralBus_oe && !peripheralBus_we;

	always @(posedge clk) begin
		if (rst) begin
			registerValue <= DEFAULT;
		end else begin
			if (we) begin
				if (enableWrite) registerValue <= writeData[WIDTH-1:0];
				else if (enableSet) registerValue <= setData;
				else if (enableClear) registerValue <= clearData;
				else if (enableToggle) registerValue <= toggleData;
			end
		end
	end

	wire[31:0] baseReadData;
	generate
		if (WIDTH == 32) begin
			assign baseReadData = registerValue;
		end else begin
			wire[32-WIDTH-1:0] zeroPadding = 'b0;
			assign baseReadData = { zeroPadding, registerValue };
		end
	endgenerate

	assign peripheralBus_dataRead = oe ? baseReadData & dataMask : 32'b0;
	assign requestOutput = oe;
	assign currentValue = registerValue;

endmodulemodule DeviceSelect #(
		parameter ID = 4'h0
	)(
		input wire peripheralEnable,
		input wire[15:0] peripheralBus_address,
		output wire[11:0] localAddress,
		output wire deviceEnable
	);

	assign deviceEnable = peripheralEnable && (peripheralBus_address[15:12] == ID);
	assign localAddress = peripheralBus_address[11:0];

endmodulemodule PeripheralSelect #(
		parameter ID = 8'h00
	)(
		input wire[23:0] peripheralBus_address,
		output wire[15:0] localAddress,
		output wire peripheralEnable
	);

	assign peripheralEnable = peripheralBus_address[23:16] == ID;
	assign localAddress = peripheralBus_address[15:0];

endmodulemodule Video (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground

		input wire wb_clk_i,
		input wire wb_rst_i,

		// Wishbone Slave ports
		input wire wb_stb_i,
		input wire wb_cyc_i,
		input wire wb_we_i,
		input wire[3:0] wb_sel_i,
		input wire[31:0] wb_data_i,
		input wire[23:0] wb_adr_i,
		output wire wb_ack_o,
		output wire wb_stall_o,
		output wire wb_error_o,
		output wire[31:0] wb_data_o,

		// IRQ
		output wire[1:0] video_irq,

		// Left Video SRAM rw port
		output wire sram0_clk0,
		output wire[1:0] sram0_csb0,
		output wire sram0_web0,
		output wire[3:0] sram0_wmask0,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram0_addr0,
		output wire[31:0] sram0_din0,
		input wire[63:0] sram0_dout0,

		// Left Video SRAM r port
		output wire sram0_clk1,
		output wire[1:0] sram0_csb1,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram0_addr1,
		input wire[63:0] sram0_dout1,

		// Right Video SRAM rw port
		output wire sram1_clk0,
		output wire[1:0] sram1_csb0,
		output wire sram1_web0,
		output wire[3:0] sram1_wmask0,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram1_addr0,
		output wire[31:0] sram1_din0,
		input wire[63:0] sram1_dout0,

		// Right Video SRAM r port
		output wire sram1_clk1,
		output wire[1:0] sram1_csb1,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram1_addr1,
		input wire[63:0] sram1_dout1,

		// VGA
		//input wire vga_clk,
		output wire[1:0] vga_r,
		output wire[1:0] vga_g,
		output wire[1:0] vga_b,
		output wire vga_vsync,
		output wire vga_hsync
	);

	localparam SRAM_ADDRESS_SIZE = 9;

	wire vga_clk = wb_clk_i;

	wire peripheralBus_we;
	wire peripheralBus_oe;
	wire peripheralBus_busy;
	wire[23:0] peripheralBus_address;
	wire[3:0] peripheralBus_byteSelect;
	wire[31:0] peripheralBus_dataRead;
	wire[31:0] peripheralBus_dataWrite;

	WBPeripheralBusInterface wbPeripheralBusInterface(
	
		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground
	
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.wb_stb_i(wb_stb_i),
		.wb_cyc_i(wb_cyc_i),
		.wb_we_i(wb_we_i),
		.wb_sel_i(wb_sel_i),
		.wb_data_i(wb_data_i),
		.wb_adr_i(wb_adr_i),
		.wb_ack_o(wb_ack_o),
		.wb_stall_o(wb_stall_o),
		.wb_error_o(wb_error_o),
		.wb_data_o(wb_data_o),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(peripheralBus_busy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(peripheralBus_dataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite));
	
	wire video_fetchData;
	wire[SRAM_ADDRESS_SIZE+3:0] vga_address;
	wire[31:0] vga_data;

	wire videoMemoryBusBusy;
	wire[31:0] videoMemoryDataRead;
	wire videoMemoryRequestOutput;
	wire vga_fetchData;
	VideoMemory videoMemory(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(videoMemoryBusBusy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(videoMemoryDataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.requestOutput(videoMemoryRequestOutput),
		.video_fetchData(vga_fetchData),
		.video_address(vga_address),
		.video_data(vga_data),
		.sram0_csb0(sram0_csb0),
		.sram0_web0(sram0_web0),
		.sram0_wmask0(sram0_wmask0),
		.sram0_addr0(sram0_addr0),
		.sram0_din0(sram0_din0),
		.sram0_dout0(sram0_dout0),
		.sram0_csb1(sram0_csb1),
		.sram0_addr1(sram0_addr1),
		.sram0_dout1(sram0_dout1),
		.sram1_csb0(sram1_csb0),
		.sram1_web0(sram1_web0),
		.sram1_wmask0(sram1_wmask0),
		.sram1_addr0(sram1_addr0),
		.sram1_din0(sram1_din0),
		.sram1_dout0(sram1_dout0),
		.sram1_csb1(sram1_csb1),
		.sram1_addr1(sram1_addr1),
		.sram1_dout1(sram1_dout1));

	assign sram0_clk0 = vga_clk;
	assign sram0_clk1 = vga_clk;
	assign sram1_clk0 = vga_clk;
	assign sram1_clk1 = vga_clk;

	wire vgaBusBusy;
	wire[31:0] vgaDataRead;
	wire vgaRequestOutput;
	VGA #(.ADDRESS_BITS(SRAM_ADDRESS_SIZE + 4)) vga(

		.vccd1(vccd1),	// User area 1 1.8V power
		.vssd1(vssd1),	// User area 1 digital ground

		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(vgaBusBusy),
		.peripheralBus_address(peripheralBus_address),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataRead(vgaDataRead),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.requestOutput(vgaRequestOutput),
		.vga_clk(vga_clk),
		.vga_fetchData(vga_fetchData),
		.vga_address(vga_address),
		.vga_data(vga_data),
		.vga_r(vga_r),
		.vga_g(vga_g),
		.vga_b(vga_b),
		.vga_vsync(vga_vsync),
		.vga_hsync(vga_hsync),
		.vga_irq(video_irq));

	assign peripheralBus_busy = videoMemoryBusBusy || vgaBusBusy;
	assign peripheralBus_dataRead = videoMemoryRequestOutput ? videoMemoryDataRead : 
									vgaRequestOutput ? vgaDataRead : ~32'b0;

endmodulemodule VideoMemory (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground

		input wire clk,
		input wire rst,

		// Peripheral bus interface
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[23:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		input wire[31:0] peripheralBus_dataWrite,
		output wire[31:0] peripheralBus_dataRead,
		output wire requestOutput,

		// Video interface
		input wire video_fetchData,
		input wire[SRAM_ADDRESS_SIZE+3:0] video_address,
		output reg[31:0] video_data,

		// Left Video SRAM rw port
		output wire[1:0] sram0_csb0,
		output wire sram0_web0,
		output wire[3:0] sram0_wmask0,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram0_addr0,
		output wire[31:0] sram0_din0,
		input wire[63:0] sram0_dout0,

		// Left Video SRAM r port
		output wire[1:0] sram0_csb1,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram0_addr1,
		input wire[63:0] sram0_dout1,

		// Right Video SRAM rw port
		output wire[1:0] sram1_csb0,
		output wire sram1_web0,
		output wire[3:0] sram1_wmask0,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram1_addr0,
		output wire[31:0] sram1_din0,
		input wire[63:0] sram1_dout0,

		// Right Video SRAM r port
		output wire[1:0] sram1_csb1,
		output wire[SRAM_ADDRESS_SIZE-1:0] sram1_addr1,
		input wire[63:0] sram1_dout1
	);

	localparam SRAM_ADDRESS_SIZE = 9;

	localparam SRAM_PERIPHERAL_BUS_ADDRESS = 11'h000;

	// Merge two ports into one
	reg[3:0] sram_csb0;
	wire sram_web0;
	wire[3:0] sram_wmask0;
	wire[SRAM_ADDRESS_SIZE-1:0] sram_addr0;
	wire[31:0] sram_din0;
	wire[127:0] sram_dout0;
	reg[3:0] sram_csb1;
	wire[SRAM_ADDRESS_SIZE-1:0] sram_addr1;
	wire[127:0] sram_dout1;

	assign sram0_csb0 = sram_csb0[1:0];
	assign sram0_web0 = sram_web0;
	assign sram0_wmask0 = sram_wmask0;
	assign sram0_addr0 = sram_addr0;
	assign sram0_din0 = sram_din0;
	assign sram0_csb1 = sram_csb1[1:0];
	assign sram0_addr1 = sram_addr1;
	assign sram1_csb0 = sram_csb0[3:2];
	assign sram1_web0 = sram_web0;
	assign sram1_wmask0 = sram_wmask0;
	assign sram1_addr0 = sram_addr0;
	assign sram1_din0 = sram_din0;
	assign sram1_csb1 = sram_csb1[3:2];
	assign sram1_addr1 = sram_addr1;

	assign sram_dout0 = { sram1_dout0, sram0_dout0 };
	assign sram_dout1 = { sram1_dout1, sram0_dout1 };

	wire peripheralBusValidAddress = peripheralBus_address[23:SRAM_ADDRESS_SIZE+4] == SRAM_PERIPHERAL_BUS_ADDRESS;
	wire peripheralBusReadEnable = peripheralBus_oe && peripheralBusValidAddress;
	wire peripheralBusWriteEnable = peripheralBus_we && peripheralBusValidAddress;
	wire peripheralBusEnableSRAM = peripheralBusReadEnable || peripheralBusWriteEnable;
	wire[1:0] peripheralBusSRAMBank = peripheralBus_address[SRAM_ADDRESS_SIZE+3:SRAM_ADDRESS_SIZE+2];

	// Set enable bit for peripheral bus port (active low)
	always @(*) begin
		if (peripheralBusEnableSRAM) begin
			case (peripheralBusSRAMBank)
				2'b00: sram_csb0 <= 4'b1110;
				2'b01: sram_csb0 <= 4'b1101;
				2'b10: sram_csb0 <= 4'b1011;
				2'b11: sram_csb0 <= 4'b0111;
			endcase
		end else begin
			sram_csb0 <= 4'b1111;
		end
	end

	// Read data only valid the clock cycle after the address is sent
	reg wbReadReady = 1'b0;
	always @(posedge clk) begin
		if (rst) wbReadReady <= 1'b0;
		else if (peripheralBusReadEnable) wbReadReady <= 1'b1;
		else wbReadReady <= 1'b0;
	end

	reg[31:0] readData;
	assign peripheralBus_dataRead = {
		peripheralBus_byteSelect[3] && wbReadReady ? readData[31:24] : 8'h00,
		peripheralBus_byteSelect[2] && wbReadReady ? readData[23:16] : 8'h00,
		peripheralBus_byteSelect[1] && wbReadReady ? readData[15:8]  : 8'h00,
		peripheralBus_byteSelect[0] && wbReadReady ? readData[7:0]   : 8'h00
	};

	assign peripheralBus_busy = peripheralBusReadEnable && !wbReadReady;
	assign requestOutput = peripheralBusReadEnable;

	assign sram_web0 	= !peripheralBusWriteEnable;
	assign sram_wmask0 	= peripheralBus_byteSelect;
	assign sram_addr0 	= peripheralBus_address[SRAM_ADDRESS_SIZE+1:2];
	assign sram_din0 	= peripheralBus_dataWrite;

	// Select return data for peripheral bus port
	always @(*) begin
		if (peripheralBusReadEnable) begin
			case (peripheralBusSRAMBank)
				2'b00: readData <= sram_dout0[31:0];
				2'b01: readData <= sram_dout0[63:32];
				2'b10: readData <= sram_dout0[95:64];
				2'b11: readData <= sram_dout0[127:96];
			endcase
		end else begin
			readData <= ~32'b0;
		end
	end

	wire[1:0] videoSRAMBank = video_address[SRAM_ADDRESS_SIZE+3:SRAM_ADDRESS_SIZE+2];

	// Set enable bit for video port (active low)
	always @(*) begin
		if (video_fetchData) begin
			case (videoSRAMBank)
				2'b00: sram_csb1 <= 4'b1110;
				2'b01: sram_csb1 <= 4'b1101;
				2'b10: sram_csb1 <= 4'b1011;
				2'b11: sram_csb1 <= 4'b0111;
			endcase
		end else begin
			sram_csb1 <= 4'b1111;
		end
	end

	assign sram_addr1 	= video_address[SRAM_ADDRESS_SIZE+1:2];

	// Select return data for video port
	always @(*) begin
		case (videoSRAMBank)
			2'b00: video_data <= sram_dout1[31:0];
			2'b01: video_data <= sram_dout1[63:32];
			2'b10: video_data <= sram_dout1[95:64];
			2'b11: video_data <= sram_dout1[127:96];
		endcase
	end

endmodulemodule VGA #(
		parameter ADDRESS_BITS = 13
	)(

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground

		input wire clk,
		input wire rst,

		// Peripheral bus for configuration
		input wire peripheralBus_we,
		input wire peripheralBus_oe,
		output wire peripheralBus_busy,
		input wire[23:0] peripheralBus_address,
		input wire[3:0] peripheralBus_byteSelect,
		input wire[31:0] peripheralBus_dataWrite,
		output reg[31:0] peripheralBus_dataRead,
		output wire requestOutput,

		// Memory interface
		input wire vga_clk,
		output wire vga_fetchData,
		output reg[ADDRESS_BITS-1:0] vga_address,
		input wire[31:0] vga_data,

		// VGA output
		output wire[1:0] vga_r,
		output wire[1:0] vga_g,
		output wire[1:0] vga_b,
		output wire vga_vsync,
		output wire vga_hsync,

		// IRQ
		output wire[1:0] vga_irq
	);
	
	// MAX_ROW_WIDTH = 2^ROW_BITS = 64;
	// MAX_COLUMN_WIDTH = 2^COLUMN_BITS * (MAX_SUB_PIXEL_VALUE+1) = 80;

	localparam VERTICAL_BITS = 7;
	localparam HORIZONTAL_BITS = 4;
	localparam MAX_SUB_PIXEL_VALUE = 3'h4;

	localparam DRAW_MODE_RAW 	 	  	= 2'b00;
	localparam DRAW_MODE_RAW_TIGHT_MEM 	= 2'b01;
	localparam DRAW_MODE_COLOUR_PALETTE = 2'b10;
	localparam DRAW_MODE_SPRITES 	  	= 2'b11;

	localparam CONFIG_ADDRESS = 12'h800;

	wire configEnable = peripheralBus_address[23:12] == CONFIG_ADDRESS;
	wire[11:0] configRegisterAddress = peripheralBus_address[11:0];

	//  Registers
	// Configuration 	Default 0x0AA
	// b00-b03: horizontalPixelSize		Default 0xA
	// b04-b07: verticalPixelSize		Default 0xA
	// b08-b09: drawMode 				Default 0b00
	// b10: enableOutput				Default 0
	// b11: hsyncInterruptEnable		Default 0
	// b12: vsyncInterruptEnable		Default 0
	wire[12:0] configuration;
	wire[31:0] configurationRegisterOutputData;
	wire configurationRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(13), .ADDRESS(12'h000), .DEFAULT(11'h0AA)) configurationRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(configurationRegisterOutputData),
		.requestOutput(configurationRegisterOutputRequest),
		.currentValue(configuration));
	
	wire[3:0] horizontalPixelSize = configuration[3:0];
	wire[3:0] verticalPixelSize   = configuration[7:4];
	wire[1:0] drawMode 			  = configuration[9:8];
	wire enableOutput 			  = configuration[10];
	wire hsyncInterruptEnable 	  = configuration[11];
	wire vsyncInterruptEnable 	  = configuration[12];

	// Defaults are timing for 800 x 600 at 60Hz
	// http://tinyvga.com/vga-timing/800x600@60Hz
	// Horizontal visible area compare 	Default 799=0x31F
	wire[10:0] horizontalVisibleAreaCompare;
	wire[31:0] horizontalVisibleAreaCompareRegisterOutputData;
	wire horizontalVisibleAreaCompareRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(11), .ADDRESS(12'h010), .DEFAULT(11'h31F)) horizontalVisibleAreaCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(horizontalVisibleAreaCompareRegisterOutputData),
		.requestOutput(horizontalVisibleAreaCompareRegisterOutputRequest),
		.currentValue(horizontalVisibleAreaCompare));

	// Horizontal front porch compare 	Default 839=0x347
	wire[10:0] horizontalFrontPorchCompare;
	wire[31:0] horizontalFrontPorchCompareRegisterOutputData;
	wire horizontalFrontPorchCompareRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(11), .ADDRESS(12'h014), .DEFAULT(11'h347)) horizontalFrontPorchCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(horizontalFrontPorchCompareRegisterOutputData),
		.requestOutput(horizontalFrontPorchCompareRegisterOutputRequest),
		.currentValue(horizontalFrontPorchCompare));

	// Horizontal sync pulse compare 	Default 967=0x3C7
	wire[10:0] horizontalSyncPulseCompare;
	wire[31:0] horizontalSyncPulseCompareRegisterOutputData;
	wire horizontalSyncPulseCompareRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(11), .ADDRESS(12'h018), .DEFAULT(11'h3C7)) horizontalSyncPulseCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(horizontalSyncPulseCompareRegisterOutputData),
		.requestOutput(horizontalSyncPulseCompareRegisterOutputRequest),
		.currentValue(horizontalSyncPulseCompare));

	// Horizontal whole line compare 	Default 1055=0x41F
	wire[10:0] horizontalWholeLineCompare;
	wire[31:0] horizontalWholeLineCompareRegisterOutputData;
	wire horizontalWholeLineCompareRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(11), .ADDRESS(12'h01C), .DEFAULT(11'h41F)) horizontalWholeLineCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(horizontalWholeLineCompareRegisterOutputData),
		.requestOutput(horizontalWholeLineCompareRegisterOutputRequest),
		.currentValue(horizontalWholeLineCompare));

	// Vertical visible area compare 	Default 599=0x257
	wire[9:0] verticalVisibleAreaCompare;
	wire[31:0] verticalVisibleAreaCompareRegisterOutputData;
	wire verticalVisibleAreaCompareRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(10), .ADDRESS(12'h020), .DEFAULT(11'h257)) verticalVisibleAreaCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(verticalVisibleAreaCompareRegisterOutputData),
		.requestOutput(verticalVisibleAreaCompareRegisterOutputRequest),
		.currentValue(verticalVisibleAreaCompare));

	// Vertical front porch compare 	Default 600=0x258
	wire[9:0] verticalFrontPorchCompare;
	wire[31:0] verticalFrontPorchCompareRegisterOutputData;
	wire verticalFrontPorchCompareRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(10), .ADDRESS(12'h024), .DEFAULT(11'h258)) verticalFrontPorchCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(verticalFrontPorchCompareRegisterOutputData),
		.requestOutput(verticalFrontPorchCompareRegisterOutputRequest),
		.currentValue(verticalFrontPorchCompare));

	// Vertical sync pulse compare 	Default 604=0x25C
	wire[9:0] verticalSyncPulseCompare;
	wire[31:0] verticalSyncPulseCompareRegisterOutputData;
	wire verticalSyncPulseCompareRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(10), .ADDRESS(12'h028), .DEFAULT(11'h25C)) verticalSyncPulseCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(verticalSyncPulseCompareRegisterOutputData),
		.requestOutput(verticalSyncPulseCompareRegisterOutputRequest),
		.currentValue(verticalSyncPulseCompare));

	// Vertical whole line compare 	Default 627=0x273
	wire[9:0] verticalWholeLineCompare;
	wire[31:0] verticalWholeLineCompareRegisterOutputData;
	wire verticalWholeLineCompareRegisterOutputRequest;
	ConfigurationRegister #(.WIDTH(10), .ADDRESS(12'h02C), .DEFAULT(11'h273)) verticalWholeLineCompareRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(verticalWholeLineCompareRegisterOutputData),
		.requestOutput(verticalWholeLineCompareRegisterOutputRequest),
		.currentValue(verticalWholeLineCompare));

	// VGA state register
	reg[4:0] stateRegisterBuffered;
	reg inVerticalVisibleArea = 1'b1;
	reg inHorizontalVisibleArea = 1'b1;
	wire[31:0] stateRegisterOutputData;
	wire stateRegisterOutputRequest;
	wire stateReadDataEnable_nc;
	wire stateRegisterBusyBusy_nc;
	wire[4:0] stateRegisterWriteData_nc;
	wire stateRegisterWriteDataEnable_nc;
	DataRegister #(.WIDTH(5), .ADDRESS(12'h030)) stateRegister(
		.clk(clk),
		.rst(rst),
		.enable(configEnable),
		.peripheralBus_we(peripheralBus_we),
		.peripheralBus_oe(peripheralBus_oe),
		.peripheralBus_busy(stateRegisterBusyBusy_nc),
		.peripheralBus_address(configRegisterAddress),
		.peripheralBus_byteSelect(peripheralBus_byteSelect),
		.peripheralBus_dataWrite(peripheralBus_dataWrite),
		.peripheralBus_dataRead(stateRegisterOutputData),
		.requestOutput(stateRegisterOutputRequest),
		.writeData(stateRegisterWriteData_nc),
		.writeData_en(stateRegisterWriteDataEnable_nc),
		.writeData_busy(1'b0),
		.readData(stateRegisterBuffered),
		.readData_en(stateReadDataEnable_nc),
		.readData_busy(1'b0));

	always @(posedge clk) begin
		if (rst) stateRegisterBuffered <= 5'b0;
		else stateRegisterBuffered <= { inVerticalVisibleArea, inHorizontalVisibleArea, !vga_vsync, !vga_hsync, enableOutput };
	end

	assign peripheralBus_busy = 1'b0;
	assign requestOutput = configurationRegisterOutputRequest
						|| horizontalVisibleAreaCompareRegisterOutputRequest
						|| horizontalFrontPorchCompareRegisterOutputRequest
						|| horizontalSyncPulseCompareRegisterOutputRequest
						|| horizontalWholeLineCompareRegisterOutputRequest
						|| verticalVisibleAreaCompareRegisterOutputRequest
						|| verticalFrontPorchCompareRegisterOutputRequest
						|| verticalSyncPulseCompareRegisterOutputRequest
						|| verticalWholeLineCompareRegisterOutputRequest
						|| stateRegisterOutputRequest;

	always @(*) begin
		case (1'b1)
			configurationRegisterOutputRequest:
				peripheralBus_dataRead <= configurationRegisterOutputData;
			horizontalVisibleAreaCompareRegisterOutputRequest:
				peripheralBus_dataRead <= horizontalVisibleAreaCompareRegisterOutputData;
			horizontalFrontPorchCompareRegisterOutputRequest:
				peripheralBus_dataRead <= horizontalFrontPorchCompareRegisterOutputData;
			horizontalSyncPulseCompareRegisterOutputRequest:
				peripheralBus_dataRead <= horizontalSyncPulseCompareRegisterOutputData;
			horizontalWholeLineCompareRegisterOutputRequest:
				peripheralBus_dataRead <= horizontalWholeLineCompareRegisterOutputData;
			verticalVisibleAreaCompareRegisterOutputRequest:
				peripheralBus_dataRead <= verticalVisibleAreaCompareRegisterOutputData;
			verticalFrontPorchCompareRegisterOutputRequest:
				peripheralBus_dataRead <= verticalFrontPorchCompareRegisterOutputData;
			verticalSyncPulseCompareRegisterOutputRequest:
				peripheralBus_dataRead <= verticalSyncPulseCompareRegisterOutputData;
			verticalWholeLineCompareRegisterOutputRequest:
				peripheralBus_dataRead <= verticalWholeLineCompareRegisterOutputData;
			stateRegisterOutputRequest:
				peripheralBus_dataRead <= stateRegisterOutputData;
			default: peripheralBus_dataRead <= ~32'b0;
		endcase
	end

	// VGA sync signal generations
	reg[10:0] horizontalCounter;
	wire isEndHorizontalVisibleArea = horizontalCounter == horizontalVisibleAreaCompare;
	wire isEndHorizontalFrontPorch = horizontalCounter == horizontalFrontPorchCompare;
	wire isEndHorizontalSyncPulse = horizontalCounter == horizontalSyncPulseCompare;
	wire isEndHorizontalWholeLine = horizontalCounter == horizontalWholeLineCompare;

	reg hsync;
	always @(posedge vga_clk) begin
		if (rst || !enableOutput) begin
			horizontalCounter <= 10'b0;
			inHorizontalVisibleArea <= 1'b1;
			hsync <= 1'b1;
		end else begin
			if (isEndHorizontalWholeLine) horizontalCounter <= 10'b0;
			else horizontalCounter <= horizontalCounter + 1;

			if (isEndHorizontalVisibleArea) inHorizontalVisibleArea <= 1'b0;
			else if (isEndHorizontalWholeLine) inHorizontalVisibleArea <= 1'b1;

			if (isEndHorizontalFrontPorch) hsync <= 1'b0;
			else if (isEndHorizontalSyncPulse) hsync <= 1'b1;
		end
	end
	
	reg[9:0] verticalCounter;
	wire isEndVerticalVisibleArea = verticalCounter == verticalVisibleAreaCompare;
	wire isEndVerticalFrontPorch = verticalCounter == verticalFrontPorchCompare;
	wire isEndVerticalSyncPulse = verticalCounter == verticalSyncPulseCompare;
	wire isEndVerticalWholeLine = verticalCounter == verticalWholeLineCompare;

	reg vsync;
	always @(posedge vga_clk) begin
		if (rst || !enableOutput) begin
			verticalCounter <= 10'b0;
			inVerticalVisibleArea <= 1'b1;
			vsync <= 1'b1;
		end else begin
			if (isEndHorizontalWholeLine) begin
				if (isEndVerticalWholeLine) verticalCounter <= 10'b0;
				else verticalCounter <= verticalCounter + 1;

				if (isEndVerticalVisibleArea) inVerticalVisibleArea <= 1'b0;
				else if (isEndVerticalWholeLine) inVerticalVisibleArea <= 1'b1;

				if (isEndVerticalFrontPorch) vsync <= 1'b0;
				else if (isEndVerticalSyncPulse) vsync <= 1'b1;
			end
		end
	end

	// Latch data in from sram and delay sync signals
	// Data timing
	// c0: pixel counter increments, sync signal set, and address is set 
	// c1: data is valid

	reg fetchPixelData;
	reg loadPixelData;

	reg[31:0] currentPixelData;
	always @(posedge vga_clk) begin
		if (rst || !enableOutput) begin
			currentPixelData <= 32'b0;
			loadPixelData <= 1'b0;
		end else begin
			loadPixelData <= fetchPixelData;
			if (loadPixelData) currentPixelData <= vga_data;
		end
	end

	assign vga_fetchData = fetchPixelData;

	assign vga_hsync = enableOutput ? hsync : 1'b1;
	assign vga_vsync = enableOutput ? vsync : 1'b1;

	// VGA pixel address select
	reg[8:0] raw_horizontalPixelCounter;
	wire[8:0] raw_nextHorizontalPixelCounter = raw_horizontalPixelCounter + 1;
	reg[9:0] raw_verticalPixelCounter;
	reg[2:0] raw_subPixelCounter;
	reg[2:0] raw_subPixelCounter_buffered;

	reg[8:0] raw_horizontalPixelCounter_d;
	reg[9:0] raw_verticalPixelCounter_d;
	reg[2:0] raw_subPixelCounter_d;

	reg[3:0] raw_horizontalPixelStretchCounter = 4'b0;
	reg[3:0] raw_horizontalPixelStretchCounter_d;
	wire[3:0] raw_nextHorizontalPixelStretchCounter = raw_horizontalPixelStretchCounter + 1;
	reg[3:0] raw_verticalPixelStretchCounter = 4'b0;
	reg[3:0] raw_verticalPixelStretchCounter_d;
	wire[3:0] raw_nextVerticalPixelStretchCounter = raw_verticalPixelStretchCounter + 1;

	reg[17:0] raw_directPixelCounterVertical;
	reg[17:0] raw_directPixelCounterVertical_d;

	wire[17:0] raw_directPixelCounter = raw_directPixelCounterVertical_d + raw_horizontalPixelCounter_d;

	wire raw_horizontalPixelStretchNextPixel = raw_nextHorizontalPixelStretchCounter == horizontalPixelSize;
	wire raw_verticalPixelStretchNextPixel = raw_nextVerticalPixelStretchCounter == verticalPixelSize;

	// Raw draw mode
	always @(*) begin
		raw_directPixelCounterVertical_d = raw_directPixelCounterVertical;
		raw_subPixelCounter_d = raw_subPixelCounter;
		raw_horizontalPixelCounter_d = raw_horizontalPixelCounter;
		raw_horizontalPixelStretchCounter_d = raw_horizontalPixelStretchCounter;
		raw_verticalPixelCounter_d = raw_verticalPixelCounter;
		raw_verticalPixelStretchCounter_d = raw_verticalPixelStretchCounter;

		if (rst || !enableOutput || !inVerticalVisibleArea) begin
			raw_directPixelCounterVertical_d = 18'b0;		
			raw_subPixelCounter_d = 3'b0;
			raw_horizontalPixelCounter_d = 9'b0;
			raw_horizontalPixelStretchCounter_d = 4'b0;
			raw_verticalPixelCounter_d = 10'b0;
			raw_verticalPixelStretchCounter_d = 4'b0;	
		end else begin
			if (inHorizontalVisibleArea) begin
				if (raw_horizontalPixelStretchNextPixel) begin
					if (raw_subPixelCounter == MAX_SUB_PIXEL_VALUE) begin
						raw_subPixelCounter_d = 3'b0;
						raw_horizontalPixelCounter_d = raw_nextHorizontalPixelCounter;
					end	else begin
						raw_subPixelCounter_d = raw_subPixelCounter + 1;
					end

					raw_horizontalPixelStretchCounter_d = 4'b0;
				end else begin
					raw_horizontalPixelStretchCounter_d = raw_nextHorizontalPixelStretchCounter;
				end
			end else begin
				raw_subPixelCounter_d = 3'b0;
				raw_horizontalPixelCounter_d = 9'b0;
				raw_horizontalPixelStretchCounter_d = 4'b0;
			end

			if (isEndHorizontalVisibleArea) begin
				if (raw_verticalPixelStretchNextPixel) begin
					raw_directPixelCounterVertical_d = raw_directPixelCounterVertical + raw_nextHorizontalPixelCounter;
					raw_verticalPixelCounter_d = raw_verticalPixelCounter + 1;
					raw_verticalPixelStretchCounter_d = 4'b0;
				end else begin
					raw_verticalPixelStretchCounter_d = raw_nextVerticalPixelStretchCounter;
				end
			end
		end
	end

	always @(posedge vga_clk) begin
		if (rst || !enableOutput) begin
			raw_directPixelCounterVertical <= 18'b0;
			raw_horizontalPixelCounter <= 9'b0;
			raw_verticalPixelCounter <= 10'b0;
			raw_subPixelCounter <= 3'b0;
			raw_horizontalPixelStretchCounter <= 4'b0;
			raw_verticalPixelStretchCounter <= 4'b0;
		end else begin
			raw_directPixelCounterVertical <= raw_directPixelCounterVertical_d;
			raw_horizontalPixelCounter <= raw_horizontalPixelCounter_d;
			raw_verticalPixelCounter <= raw_verticalPixelCounter_d;
			raw_subPixelCounter <= raw_subPixelCounter_d;
			raw_subPixelCounter_buffered <= raw_subPixelCounter;
			raw_horizontalPixelStretchCounter <= raw_horizontalPixelStretchCounter_d;
			raw_verticalPixelStretchCounter <= raw_verticalPixelStretchCounter_d;
		end
	end

	wire raw_verticalPixelCounterChanged = raw_verticalPixelCounter != raw_verticalPixelCounter_d;
	wire raw_horizontalPixelCounterChanged = raw_horizontalPixelCounter != raw_horizontalPixelCounter_d;
	wire raw_directPixelCounterChanged = raw_verticalPixelCounterChanged || raw_horizontalPixelCounterChanged;

	always @(*) begin
		if (rst || !enableOutput) begin
			vga_address <= {ADDRESS_BITS{1'b0}};
			fetchPixelData <= 1'b0;
		end else begin
			// Use data register inputs for new address
			// This means that the address gets updated at the same time as the pixel counters
			// And so the data is valid the cycle after
			// Rather than being two cycles after
			case (drawMode)
				// Use Seperate horizontal and vertical portions of address
				// This means that for some resolutions portions of memory are not used by the video device
				DRAW_MODE_RAW: begin
					vga_address <= { raw_verticalPixelCounter_d[VERTICAL_BITS-1:0], raw_horizontalPixelCounter_d[HORIZONTAL_BITS-1:0], 2'b00 };
					fetchPixelData <= raw_verticalPixelCounterChanged || raw_horizontalPixelCounterChanged;
				end

				// Directly use the pixel index to access memory
				// This better uses memory, but is also slightly more complex for the cpu to write to the frame buffer
				DRAW_MODE_RAW_TIGHT_MEM: begin
					vga_address <= { raw_directPixelCounter[ADDRESS_BITS-1:0], 2'b00 };
					fetchPixelData <= raw_directPixelCounterChanged;
				end

				// TODO: Use some portion of memory to store colours, then index them with the frame buffer
				// This will require loading the pixel information ahead of time, so that the correct colour can be found
				// Is this really helpful, as we use 6-bit colour, so probably need to use 4-bit colour palette index
				DRAW_MODE_COLOUR_PALETTE: begin
					vga_address <= { raw_verticalPixelCounter_d[VERTICAL_BITS-1:0], raw_horizontalPixelCounter_d[HORIZONTAL_BITS-1:0], 2'b00 };
					fetchPixelData <= raw_verticalPixelCounterChanged || raw_horizontalPixelCounterChanged;
				end

				// TODO: Use some portion of memory to store sprites
				// Then use a sprite index rather than colour data or a colour index
				// How many sprites do we want to allow
				// How big will sprites be
				// How configurable should this be
				// We have very little video memory, so this may not work very well at all
				DRAW_MODE_SPRITES: begin
					vga_address <= { raw_verticalPixelCounter_d[VERTICAL_BITS-1:0], raw_horizontalPixelCounter_d[HORIZONTAL_BITS-1:0], 2'b00 };
					fetchPixelData <= raw_verticalPixelCounterChanged || raw_horizontalPixelCounterChanged;
				end

				default: begin
					vga_address <= { raw_verticalPixelCounter_d[VERTICAL_BITS-1:0], raw_horizontalPixelCounter_d[HORIZONTAL_BITS-1:0], 2'b00 };
					fetchPixelData <= raw_verticalPixelCounterChanged || raw_horizontalPixelCounterChanged;
				end
			endcase
		end
	end

	reg[5:0] raw_currentPixel;	
	always @(*) begin
		case (raw_subPixelCounter_buffered)
			4'h0: raw_currentPixel <= currentPixelData[5:0];
			4'h1: raw_currentPixel <= currentPixelData[11:6];
			4'h2: raw_currentPixel <= currentPixelData[17:12];
			4'h3: raw_currentPixel <= currentPixelData[23:18];
			4'h4: raw_currentPixel <= currentPixelData[29:24];
			default: raw_currentPixel <= currentPixelData[5:0];
		endcase
	end

	wire onScreen = inHorizontalVisibleArea && inVerticalVisibleArea;

	assign vga_r = enableOutput && onScreen ? raw_currentPixel[1:0] : 2'b0;
	assign vga_g = enableOutput && onScreen ? raw_currentPixel[3:2] : 2'b0;
	assign vga_b = enableOutput && onScreen ? raw_currentPixel[5:4] : 2'b0;

	// IRQ
	reg lastVSync;
	reg lastHSync;
	always @(posedge clk) begin
		if (rst) begin
			lastVSync <= 1'b0;
			lastHSync <= 1'b0;
		end else begin
			lastVSync <= vsync;
			lastHSync <= hsync;
		end
	end

	wire vsync_irq = (lastVSync != vsync) && !vsync;
	wire hsync_irq = (lastHSync != hsync) && !hsync;
	assign vga_irq = { vsync_irq && vsyncInterruptEnable, hsync_irq && hsyncInterruptEnable };

endmodule
module WishboneInterconnect (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1,	// User area 1 digital ground


		input wire wb_clk_i,
		input wire wb_rst_i,

		// Master 0
		input wire master0_wb_cyc_o,
		input wire master0_wb_stb_o,
		input wire master0_wb_we_o,
		input wire[3:0] master0_wb_sel_o,
		input wire[31:0] master0_wb_data_o,
		input wire[27:0] master0_wb_adr_o,
		output reg master0_wb_ack_i,
		output reg master0_wb_stall_i,
		output reg master0_wb_error_i,
		output reg[31:0] master0_wb_data_i,

		// Master 1
		input wire master1_wb_cyc_o,
		input wire master1_wb_stb_o,
		input wire master1_wb_we_o,
		input wire[3:0] master1_wb_sel_o,
		input wire[31:0] master1_wb_data_o,
		input wire[27:0] master1_wb_adr_o,
		output reg master1_wb_ack_i,
		output reg master1_wb_stall_i,
		output reg master1_wb_error_i,
		output reg[31:0] master1_wb_data_i,

		// Master 2
		input wire master2_wb_cyc_o,
		input wire master2_wb_stb_o,
		input wire master2_wb_we_o,
		input wire[3:0] master2_wb_sel_o,
		input wire[31:0] master2_wb_data_o,
		input wire[27:0] master2_wb_adr_o,
		output reg master2_wb_ack_i,
		output reg master2_wb_stall_i,
		output reg master2_wb_error_i,
		output reg[31:0] master2_wb_data_i,

		// Master 3
		// input wire master3_wb_cyc_o,
		// input wire master3_wb_stb_o,
		// input wire master3_wb_we_o,
		// input wire[3:0] master3_wb_sel_o,
		// input wire[31:0] master3_wb_data_o,
		// input wire[27:0] master3_wb_adr_o,
		// output reg master3_wb_ack_i,
		// output reg master3_wb_stall_i,
		// output reg master3_wb_error_i,
		// output reg[31:0] master3_wb_data_i,

		// Slave 0
		output wire slave0_wb_cyc_i,
		output wire slave0_wb_stb_i,
		output wire slave0_wb_we_i,
		output wire[3:0] slave0_wb_sel_i,
		output wire[31:0] slave0_wb_data_i,
		output wire[23:0] slave0_wb_adr_i,
		input wire slave0_wb_ack_o,
		input wire slave0_wb_stall_o,
		input wire slave0_wb_error_o,
		input wire[31:0] slave0_wb_data_o,

		// Slave 1
		output wire slave1_wb_cyc_i,
		output wire slave1_wb_stb_i,
		output wire slave1_wb_we_i,
		output wire[3:0] slave1_wb_sel_i,
		output wire[31:0] slave1_wb_data_i,
		output wire[23:0] slave1_wb_adr_i,
		input wire slave1_wb_ack_o,
		input wire slave1_wb_stall_o,
		input wire slave1_wb_error_o,
		input wire[31:0] slave1_wb_data_o,

		// Slave 2
		output wire slave2_wb_cyc_i,
		output wire slave2_wb_stb_i,
		output wire slave2_wb_we_i,
		output wire[3:0] slave2_wb_sel_i,
		output wire[31:0] slave2_wb_data_i,
		output wire[23:0] slave2_wb_adr_i,
		input wire slave2_wb_ack_o,
		input wire slave2_wb_stall_o,
		input wire slave2_wb_error_o,
		input wire[31:0] slave2_wb_data_o,

		// Slave 3
		output wire slave3_wb_cyc_i,
		output wire slave3_wb_stb_i,
		output wire slave3_wb_we_i,
		output wire[3:0] slave3_wb_sel_i,
		output wire[31:0] slave3_wb_data_i,
		output wire[23:0] slave3_wb_adr_i,
		input wire slave3_wb_ack_o,
		input wire slave3_wb_stall_o,
		input wire slave3_wb_error_o,
		input wire[31:0] slave3_wb_data_o,

		// Slave 4
		output wire slave4_wb_cyc_i,
		output wire slave4_wb_stb_i,
		output wire slave4_wb_we_i,
		output wire[3:0] slave4_wb_sel_i,
		output wire[31:0] slave4_wb_data_i,
		output wire[23:0] slave4_wb_adr_i,
		input wire slave4_wb_ack_o,
		input wire slave4_wb_stall_o,
		input wire slave4_wb_error_o,
		input wire[31:0] slave4_wb_data_o,

		// output wire[2:0] probe_master0_currentSlave,
		// output wire[2:0] probe_master1_currentSlave,
		// output wire[2:0] probe_master2_currentSlave,
		// output wire[2:0] probe_master3_currentSlave,
		// output wire[1:0] probe_slave0_currentMaster,
		// output wire[1:0] probe_slave1_currentMaster,
		// output wire[1:0] probe_slave2_currentMaster,
		// output wire[1:0] probe_slave3_currentMaster,
		// output wire[1:0] probe_slave4_currentMaster
		output wire[1:0] probe_master0_currentSlave,
		output wire[1:0] probe_master1_currentSlave,
		output wire[1:0] probe_master2_currentSlave,
		output wire[1:0] probe_master3_currentSlave,
		output wire[1:0] probe_slave0_currentMaster,
		output wire[1:0] probe_slave1_currentMaster,
		output wire[1:0] probe_slave2_currentMaster,
		output wire[1:0] probe_slave3_currentMaster
	);

	localparam SLAVE0_ADDRESS = 4'h0;
	localparam SLAVE1_ADDRESS = 4'h1;
	localparam SLAVE2_ADDRESS = 4'h2;
	localparam SLAVE3_ADDRESS = 4'h3;
	localparam SLAVE4_ADDRESS = 4'h4;

	// Disble master3
	wire master3_wb_cyc_o = 1'b0;
	wire master3_wb_stb_o = 1'b0;
	wire master3_wb_we_o = 1'b0;
	wire[3:0] master3_wb_sel_o = 4'b0;
	wire[31:0] master3_wb_data_o = ~32'b0;
	wire[27:0] master3_wb_adr_o = 28'b0;
	reg master3_wb_ack_i;
	reg master3_wb_stall_i;
	reg master3_wb_error_i;
	reg[31:0] master3_wb_data_i;

	// Master select signals
	// Master 0
	wire master0_slave0_select = master0_wb_adr_o[27:24] == SLAVE0_ADDRESS;
	wire master0_slave1_select = master0_wb_adr_o[27:24] == SLAVE1_ADDRESS;
	wire master0_slave2_select = master0_wb_adr_o[27:24] == SLAVE2_ADDRESS;
	wire master0_slave3_select = master0_wb_adr_o[27:24] == SLAVE3_ADDRESS;
	wire master0_slave4_select = master0_wb_adr_o[27:24] == SLAVE4_ADDRESS;

	// Master 1
	wire master1_slave0_select = master1_wb_adr_o[27:24] == SLAVE0_ADDRESS;
	wire master1_slave1_select = master1_wb_adr_o[27:24] == SLAVE1_ADDRESS;
	wire master1_slave2_select = master1_wb_adr_o[27:24] == SLAVE2_ADDRESS;
	wire master1_slave3_select = master1_wb_adr_o[27:24] == SLAVE3_ADDRESS;
	wire master1_slave4_select = master1_wb_adr_o[27:24] == SLAVE4_ADDRESS;

	// Master 2
	wire master2_slave0_select = master2_wb_adr_o[27:24] == SLAVE0_ADDRESS;
	wire master2_slave1_select = master2_wb_adr_o[27:24] == SLAVE1_ADDRESS;
	wire master2_slave2_select = master2_wb_adr_o[27:24] == SLAVE2_ADDRESS;
	wire master2_slave3_select = master2_wb_adr_o[27:24] == SLAVE3_ADDRESS;
	wire master2_slave4_select = master2_wb_adr_o[27:24] == SLAVE4_ADDRESS;

	// Master 3
	wire master3_slave0_select = master3_wb_adr_o[27:24] == SLAVE0_ADDRESS;
	wire master3_slave1_select = master3_wb_adr_o[27:24] == SLAVE1_ADDRESS;
	wire master3_slave2_select = master3_wb_adr_o[27:24] == SLAVE2_ADDRESS;
	wire master3_slave3_select = master3_wb_adr_o[27:24] == SLAVE3_ADDRESS;
	wire master3_slave4_select = master3_wb_adr_o[27:24] == SLAVE4_ADDRESS;

	// Slave return signals
	// Master 0
	wire master0_slave0_wb_ack_i;
	wire master0_slave0_wb_stall_i;
	wire master0_slave0_wb_error_i;
	wire[31:0] master0_slave0_wb_data_i;
	wire master0_slave1_wb_ack_i;
	wire master0_slave1_wb_stall_i;
	wire master0_slave1_wb_error_i;
	wire[31:0] master0_slave1_wb_data_i;
	wire master0_slave2_wb_ack_i;
	wire master0_slave2_wb_stall_i;
	wire master0_slave2_wb_error_i;
	wire[31:0] master0_slave2_wb_data_i;
	wire master0_slave3_wb_ack_i;
	wire master0_slave3_wb_stall_i;
	wire master0_slave3_wb_error_i;
	wire[31:0] master0_slave3_wb_data_i;
	wire master0_slave4_wb_ack_i;
	wire master0_slave4_wb_stall_i;
	wire master0_slave4_wb_error_i;
	wire[31:0] master0_slave4_wb_data_i;

	// Master 1
	wire master1_slave0_wb_ack_i;
	wire master1_slave0_wb_stall_i;
	wire master1_slave0_wb_error_i;
	wire[31:0] master1_slave0_wb_data_i;
	wire master1_slave1_wb_ack_i;
	wire master1_slave1_wb_stall_i;
	wire master1_slave1_wb_error_i;
	wire[31:0] master1_slave1_wb_data_i;
	wire master1_slave2_wb_ack_i;
	wire master1_slave2_wb_stall_i;
	wire master1_slave2_wb_error_i;
	wire[31:0] master1_slave2_wb_data_i;
	wire master1_slave3_wb_ack_i;
	wire master1_slave3_wb_stall_i;
	wire master1_slave3_wb_error_i;
	wire[31:0] master1_slave3_wb_data_i;
	wire master1_slave4_wb_ack_i;
	wire master1_slave4_wb_stall_i;
	wire master1_slave4_wb_error_i;
	wire[31:0] master1_slave4_wb_data_i;

	// Master 2
	wire master2_slave0_wb_ack_i;
	wire master2_slave0_wb_stall_i;
	wire master2_slave0_wb_error_i;
	wire[31:0] master2_slave0_wb_data_i;
	wire master2_slave1_wb_ack_i;
	wire master2_slave1_wb_stall_i;
	wire master2_slave1_wb_error_i;
	wire[31:0] master2_slave1_wb_data_i;
	wire master2_slave2_wb_ack_i;
	wire master2_slave2_wb_stall_i;
	wire master2_slave2_wb_error_i;
	wire[31:0] master2_slave2_wb_data_i;
	wire master2_slave3_wb_ack_i;
	wire master2_slave3_wb_stall_i;
	wire master2_slave3_wb_error_i;
	wire[31:0] master2_slave3_wb_data_i;
	wire master2_slave4_wb_ack_i;
	wire master2_slave4_wb_stall_i;
	wire master2_slave4_wb_error_i;
	wire[31:0] master2_slave4_wb_data_i;

	// Master 3
	wire master3_slave0_wb_ack_i;
	wire master3_slave0_wb_stall_i;
	wire master3_slave0_wb_error_i;
	wire[31:0] master3_slave0_wb_data_i;
	wire master3_slave1_wb_ack_i;
	wire master3_slave1_wb_stall_i;
	wire master3_slave1_wb_error_i;
	wire[31:0] master3_slave1_wb_data_i;
	wire master3_slave2_wb_ack_i;
	wire master3_slave2_wb_stall_i;
	wire master3_slave2_wb_error_i;
	wire[31:0] master3_slave2_wb_data_i;
	wire master3_slave3_wb_ack_i;
	wire master3_slave3_wb_stall_i;
	wire master3_slave3_wb_error_i;
	wire[31:0] master3_slave3_wb_data_i;
	wire master3_slave4_wb_ack_i;
	wire master3_slave4_wb_stall_i;
	wire master3_slave4_wb_error_i;
	wire[31:0] master3_slave4_wb_data_i;

	// Slave 0
	WishboneMultiMasterSlave slave0MultiMaster(
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.master0_wb_cyc_o(master0_wb_cyc_o && master0_slave0_select),
		.master0_wb_stb_o(master0_wb_stb_o),
		.master0_wb_we_o(master0_wb_we_o),
		.master0_wb_sel_o(master0_wb_sel_o),
		.master0_wb_data_o(master0_wb_data_o),
		.master0_wb_adr_o(master0_wb_adr_o[23:0]),
		.master0_wb_ack_i(master0_slave0_wb_ack_i),
		.master0_wb_stall_i(master0_slave0_wb_stall_i),
		.master0_wb_error_i(master0_slave0_wb_error_i),
		.master0_wb_data_i(master0_slave0_wb_data_i),
		.master1_wb_cyc_o(master1_wb_cyc_o && master1_slave0_select),
		.master1_wb_stb_o(master1_wb_stb_o),
		.master1_wb_we_o(master1_wb_we_o),
		.master1_wb_sel_o(master1_wb_sel_o),
		.master1_wb_data_o(master1_wb_data_o),
		.master1_wb_adr_o(master1_wb_adr_o[23:0]),
		.master1_wb_ack_i(master1_slave0_wb_ack_i),
		.master1_wb_stall_i(master1_slave0_wb_stall_i),
		.master1_wb_error_i(master1_slave0_wb_error_i),
		.master1_wb_data_i(master1_slave0_wb_data_i),
		.master2_wb_cyc_o(master2_wb_cyc_o && master2_slave0_select),
		.master2_wb_stb_o(master2_wb_stb_o),
		.master2_wb_we_o(master2_wb_we_o),
		.master2_wb_sel_o(master2_wb_sel_o),
		.master2_wb_data_o(master2_wb_data_o),
		.master2_wb_adr_o(master2_wb_adr_o[23:0]),
		.master2_wb_ack_i(master2_slave0_wb_ack_i),
		.master2_wb_stall_i(master2_slave0_wb_stall_i),
		.master2_wb_error_i(master2_slave0_wb_error_i),
		.master2_wb_data_i(master2_slave0_wb_data_i),
		.master3_wb_cyc_o(master3_wb_cyc_o && master3_slave0_select),
		.master3_wb_stb_o(master3_wb_stb_o),
		.master3_wb_we_o(master3_wb_we_o),
		.master3_wb_sel_o(master3_wb_sel_o),
		.master3_wb_data_o(master3_wb_data_o),
		.master3_wb_adr_o(master3_wb_adr_o[23:0]),
		.master3_wb_ack_i(master3_slave0_wb_ack_i),
		.master3_wb_stall_i(master3_slave0_wb_stall_i),
		.master3_wb_error_i(master3_slave0_wb_error_i),
		.master3_wb_data_i(master3_slave0_wb_data_i),
		.slave_cyc_i(slave0_wb_cyc_i),
		.slave_stb_i(slave0_wb_stb_i),
		.slave_we_i(slave0_wb_we_i),
		.slave_sel_i(slave0_wb_sel_i),
		.slave_data_i(slave0_wb_data_i),
		.slave_adr_i(slave0_wb_adr_i),
		.slave_ack_o(slave0_wb_ack_o),
		.slave_stall_o(slave0_wb_stall_o),
		.slave_error_o(slave0_wb_error_o),
		.slave_data_o(slave0_wb_data_o),
		.probe_currentMaster(probe_slave0_currentMaster));

	// Slave 1
	WishboneMultiMasterSlave slave1MultiMaster(
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.master0_wb_cyc_o(master0_wb_cyc_o && master0_slave1_select),
		.master0_wb_stb_o(master0_wb_stb_o),
		.master0_wb_we_o(master0_wb_we_o),
		.master0_wb_sel_o(master0_wb_sel_o),
		.master0_wb_data_o(master0_wb_data_o),
		.master0_wb_adr_o(master0_wb_adr_o[23:0]),
		.master0_wb_ack_i(master0_slave1_wb_ack_i),
		.master0_wb_stall_i(master0_slave1_wb_stall_i),
		.master0_wb_error_i(master0_slave1_wb_error_i),
		.master0_wb_data_i(master0_slave1_wb_data_i),
		.master1_wb_cyc_o(master1_wb_cyc_o && master1_slave1_select),
		.master1_wb_stb_o(master1_wb_stb_o),
		.master1_wb_we_o(master1_wb_we_o),
		.master1_wb_sel_o(master1_wb_sel_o),
		.master1_wb_data_o(master1_wb_data_o),
		.master1_wb_adr_o(master1_wb_adr_o[23:0]),
		.master1_wb_ack_i(master1_slave1_wb_ack_i),
		.master1_wb_stall_i(master1_slave1_wb_stall_i),
		.master1_wb_error_i(master1_slave1_wb_error_i),
		.master1_wb_data_i(master1_slave1_wb_data_i),
		.master2_wb_cyc_o(master2_wb_cyc_o && master2_slave1_select),
		.master2_wb_stb_o(master2_wb_stb_o),
		.master2_wb_we_o(master2_wb_we_o),
		.master2_wb_sel_o(master2_wb_sel_o),
		.master2_wb_data_o(master2_wb_data_o),
		.master2_wb_adr_o(master2_wb_adr_o[23:0]),
		.master2_wb_ack_i(master2_slave1_wb_ack_i),
		.master2_wb_stall_i(master2_slave1_wb_stall_i),
		.master2_wb_error_i(master2_slave1_wb_error_i),
		.master2_wb_data_i(master2_slave1_wb_data_i),
		.master3_wb_cyc_o(master3_wb_cyc_o && master3_slave1_select),
		.master3_wb_stb_o(master3_wb_stb_o),
		.master3_wb_we_o(master3_wb_we_o),
		.master3_wb_sel_o(master3_wb_sel_o),
		.master3_wb_data_o(master3_wb_data_o),
		.master3_wb_adr_o(master3_wb_adr_o[23:0]),
		.master3_wb_ack_i(master3_slave1_wb_ack_i),
		.master3_wb_stall_i(master3_slave1_wb_stall_i),
		.master3_wb_error_i(master3_slave1_wb_error_i),
		.master3_wb_data_i(master3_slave1_wb_data_i),
		.slave_cyc_i(slave1_wb_cyc_i),
		.slave_stb_i(slave1_wb_stb_i),
		.slave_we_i(slave1_wb_we_i),
		.slave_sel_i(slave1_wb_sel_i),
		.slave_data_i(slave1_wb_data_i),
		.slave_adr_i(slave1_wb_adr_i),
		.slave_ack_o(slave1_wb_ack_o),
		.slave_stall_o(slave1_wb_stall_o),
		.slave_error_o(slave1_wb_error_o),
		.slave_data_o(slave1_wb_data_o),
		.probe_currentMaster(probe_slave1_currentMaster));

	// Slave 2
	WishboneMultiMasterSlave slave2MultiMaster(
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.master0_wb_cyc_o(master0_wb_cyc_o && master0_slave2_select),
		.master0_wb_stb_o(master0_wb_stb_o),
		.master0_wb_we_o(master0_wb_we_o),
		.master0_wb_sel_o(master0_wb_sel_o),
		.master0_wb_data_o(master0_wb_data_o),
		.master0_wb_adr_o(master0_wb_adr_o[23:0]),
		.master0_wb_ack_i(master0_slave2_wb_ack_i),
		.master0_wb_stall_i(master0_slave2_wb_stall_i),
		.master0_wb_error_i(master0_slave2_wb_error_i),
		.master0_wb_data_i(master0_slave2_wb_data_i),
		.master1_wb_cyc_o(master1_wb_cyc_o && master1_slave2_select),
		.master1_wb_stb_o(master1_wb_stb_o),
		.master1_wb_we_o(master1_wb_we_o),
		.master1_wb_sel_o(master1_wb_sel_o),
		.master1_wb_data_o(master1_wb_data_o),
		.master1_wb_adr_o(master1_wb_adr_o[23:0]),
		.master1_wb_ack_i(master1_slave2_wb_ack_i),
		.master1_wb_stall_i(master1_slave2_wb_stall_i),
		.master1_wb_error_i(master1_slave2_wb_error_i),
		.master1_wb_data_i(master1_slave2_wb_data_i),
		.master2_wb_cyc_o(master2_wb_cyc_o && master2_slave2_select),
		.master2_wb_stb_o(master2_wb_stb_o),
		.master2_wb_we_o(master2_wb_we_o),
		.master2_wb_sel_o(master2_wb_sel_o),
		.master2_wb_data_o(master2_wb_data_o),
		.master2_wb_adr_o(master2_wb_adr_o[23:0]),
		.master2_wb_ack_i(master2_slave2_wb_ack_i),
		.master2_wb_stall_i(master2_slave2_wb_stall_i),
		.master2_wb_error_i(master2_slave2_wb_error_i),
		.master2_wb_data_i(master2_slave2_wb_data_i),
		.master3_wb_cyc_o(master3_wb_cyc_o && master3_slave2_select),
		.master3_wb_stb_o(master3_wb_stb_o),
		.master3_wb_we_o(master3_wb_we_o),
		.master3_wb_sel_o(master3_wb_sel_o),
		.master3_wb_data_o(master3_wb_data_o),
		.master3_wb_adr_o(master3_wb_adr_o[23:0]),
		.master3_wb_ack_i(master3_slave2_wb_ack_i),
		.master3_wb_stall_i(master3_slave2_wb_stall_i),
		.master3_wb_error_i(master3_slave2_wb_error_i),
		.master3_wb_data_i(master3_slave2_wb_data_i),
		.slave_cyc_i(slave2_wb_cyc_i),
		.slave_stb_i(slave2_wb_stb_i),
		.slave_we_i(slave2_wb_we_i),
		.slave_sel_i(slave2_wb_sel_i),
		.slave_data_i(slave2_wb_data_i),
		.slave_adr_i(slave2_wb_adr_i),
		.slave_ack_o(slave2_wb_ack_o),
		.slave_stall_o(slave2_wb_stall_o),
		.slave_error_o(slave2_wb_error_o),
		.slave_data_o(slave2_wb_data_o),
		.probe_currentMaster(probe_slave2_currentMaster));

	// Slave 3
	WishboneMultiMasterSlave slave3MultiMaster(
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.master0_wb_cyc_o(master0_wb_cyc_o && master0_slave3_select),
		.master0_wb_stb_o(master0_wb_stb_o),
		.master0_wb_we_o(master0_wb_we_o),
		.master0_wb_sel_o(master0_wb_sel_o),
		.master0_wb_data_o(master0_wb_data_o),
		.master0_wb_adr_o(master0_wb_adr_o[23:0]),
		.master0_wb_ack_i(master0_slave3_wb_ack_i),
		.master0_wb_stall_i(master0_slave3_wb_stall_i),
		.master0_wb_error_i(master0_slave3_wb_error_i),
		.master0_wb_data_i(master0_slave3_wb_data_i),
		.master1_wb_cyc_o(master1_wb_cyc_o && master1_slave3_select),
		.master1_wb_stb_o(master1_wb_stb_o),
		.master1_wb_we_o(master1_wb_we_o),
		.master1_wb_sel_o(master1_wb_sel_o),
		.master1_wb_data_o(master1_wb_data_o),
		.master1_wb_adr_o(master1_wb_adr_o[23:0]),
		.master1_wb_ack_i(master1_slave3_wb_ack_i),
		.master1_wb_stall_i(master1_slave3_wb_stall_i),
		.master1_wb_error_i(master1_slave3_wb_error_i),
		.master1_wb_data_i(master1_slave3_wb_data_i),
		.master2_wb_cyc_o(master2_wb_cyc_o && master2_slave3_select),
		.master2_wb_stb_o(master2_wb_stb_o),
		.master2_wb_we_o(master2_wb_we_o),
		.master2_wb_sel_o(master2_wb_sel_o),
		.master2_wb_data_o(master2_wb_data_o),
		.master2_wb_adr_o(master2_wb_adr_o[23:0]),
		.master2_wb_ack_i(master2_slave3_wb_ack_i),
		.master2_wb_stall_i(master2_slave3_wb_stall_i),
		.master2_wb_error_i(master2_slave3_wb_error_i),
		.master2_wb_data_i(master2_slave3_wb_data_i),
		.master3_wb_cyc_o(master3_wb_cyc_o && master3_slave3_select),
		.master3_wb_stb_o(master3_wb_stb_o),
		.master3_wb_we_o(master3_wb_we_o),
		.master3_wb_sel_o(master3_wb_sel_o),
		.master3_wb_data_o(master3_wb_data_o),
		.master3_wb_adr_o(master3_wb_adr_o[23:0]),
		.master3_wb_ack_i(master3_slave3_wb_ack_i),
		.master3_wb_stall_i(master3_slave3_wb_stall_i),
		.master3_wb_error_i(master3_slave3_wb_error_i),
		.master3_wb_data_i(master3_slave3_wb_data_i),
		.slave_cyc_i(slave3_wb_cyc_i),
		.slave_stb_i(slave3_wb_stb_i),
		.slave_we_i(slave3_wb_we_i),
		.slave_sel_i(slave3_wb_sel_i),
		.slave_data_i(slave3_wb_data_i),
		.slave_adr_i(slave3_wb_adr_i),
		.slave_ack_o(slave3_wb_ack_o),
		.slave_stall_o(slave3_wb_stall_o),
		.slave_error_o(slave3_wb_error_o),
		.slave_data_o(slave3_wb_data_o),
		.probe_currentMaster(probe_slave3_currentMaster));

	// Slave 4
	wire[1:0] probe_slave4_currentMaster;
	WishboneMultiMasterSlave slave4MultiMaster(
		.wb_clk_i(wb_clk_i),
		.wb_rst_i(wb_rst_i),
		.master0_wb_cyc_o(master0_wb_cyc_o && master0_slave4_select),
		.master0_wb_stb_o(master0_wb_stb_o),
		.master0_wb_we_o(master0_wb_we_o),
		.master0_wb_sel_o(master0_wb_sel_o),
		.master0_wb_data_o(master0_wb_data_o),
		.master0_wb_adr_o(master0_wb_adr_o[23:0]),
		.master0_wb_ack_i(master0_slave4_wb_ack_i),
		.master0_wb_stall_i(master0_slave4_wb_stall_i),
		.master0_wb_error_i(master0_slave4_wb_error_i),
		.master0_wb_data_i(master0_slave4_wb_data_i),
		.master1_wb_cyc_o(master1_wb_cyc_o && master1_slave4_select),
		.master1_wb_stb_o(master1_wb_stb_o),
		.master1_wb_we_o(master1_wb_we_o),
		.master1_wb_sel_o(master1_wb_sel_o),
		.master1_wb_data_o(master1_wb_data_o),
		.master1_wb_adr_o(master1_wb_adr_o[23:0]),
		.master1_wb_ack_i(master1_slave4_wb_ack_i),
		.master1_wb_stall_i(master1_slave4_wb_stall_i),
		.master1_wb_error_i(master1_slave4_wb_error_i),
		.master1_wb_data_i(master1_slave4_wb_data_i),
		.master2_wb_cyc_o(master2_wb_cyc_o && master2_slave4_select),
		.master2_wb_stb_o(master2_wb_stb_o),
		.master2_wb_we_o(master2_wb_we_o),
		.master2_wb_sel_o(master2_wb_sel_o),
		.master2_wb_data_o(master2_wb_data_o),
		.master2_wb_adr_o(master2_wb_adr_o[23:0]),
		.master2_wb_ack_i(master2_slave4_wb_ack_i),
		.master2_wb_stall_i(master2_slave4_wb_stall_i),
		.master2_wb_error_i(master2_slave4_wb_error_i),
		.master2_wb_data_i(master2_slave4_wb_data_i),
		.master3_wb_cyc_o(master3_wb_cyc_o && master3_slave4_select),
		.master3_wb_stb_o(master3_wb_stb_o),
		.master3_wb_we_o(master3_wb_we_o),
		.master3_wb_sel_o(master3_wb_sel_o),
		.master3_wb_data_o(master3_wb_data_o),
		.master3_wb_adr_o(master3_wb_adr_o[23:0]),
		.master3_wb_ack_i(master3_slave4_wb_ack_i),
		.master3_wb_stall_i(master3_slave4_wb_stall_i),
		.master3_wb_error_i(master3_slave4_wb_error_i),
		.master3_wb_data_i(master3_slave4_wb_data_i),
		.slave_cyc_i(slave4_wb_cyc_i),
		.slave_stb_i(slave4_wb_stb_i),
		.slave_we_i(slave4_wb_we_i),
		.slave_sel_i(slave4_wb_sel_i),
		.slave_data_i(slave4_wb_data_i),
		.slave_adr_i(slave4_wb_adr_i),
		.slave_ack_o(slave4_wb_ack_o),
		.slave_stall_o(slave4_wb_stall_o),
		.slave_error_o(slave4_wb_error_o),
		.slave_data_o(slave4_wb_data_o),
		.probe_currentMaster(probe_slave4_currentMaster));

	// Multiplex the connections back from the slave
	// Master 0
	always @(*) begin
		case (1'b1)
			master0_slave0_select: begin
				master0_wb_ack_i <= master0_slave0_wb_ack_i;
				master0_wb_stall_i <= master0_slave0_wb_stall_i;
				master0_wb_error_i <= master0_slave0_wb_error_i;
				master0_wb_data_i <= master0_slave0_wb_data_i;
			end
			
			master0_slave1_select: begin
				master0_wb_ack_i <= master0_slave1_wb_ack_i;
				master0_wb_stall_i <= master0_slave1_wb_stall_i;
				master0_wb_error_i <= master0_slave1_wb_error_i;
				master0_wb_data_i <= master0_slave1_wb_data_i;
			end
			
			master0_slave2_select: begin
				master0_wb_ack_i <= master0_slave2_wb_ack_i;
				master0_wb_stall_i <= master0_slave2_wb_stall_i;
				master0_wb_error_i <= master0_slave2_wb_error_i;
				master0_wb_data_i <= master0_slave2_wb_data_i;
			end
			
			master0_slave3_select: begin
				master0_wb_ack_i <= master0_slave3_wb_ack_i;
				master0_wb_stall_i <= master0_slave3_wb_stall_i;
				master0_wb_error_i <= master0_slave3_wb_error_i;
				master0_wb_data_i <= master0_slave3_wb_data_i;
			end
			
			master0_slave4_select: begin
				master0_wb_ack_i <= master0_slave4_wb_ack_i;
				master0_wb_stall_i <= master0_slave4_wb_stall_i;
				master0_wb_error_i <= master0_slave4_wb_error_i;
				master0_wb_data_i <= master0_slave4_wb_data_i;
			end
			
			default: begin
				master0_wb_ack_i <= master0_wb_cyc_o;
				master0_wb_stall_i <= 1'b0;
				master0_wb_error_i <= 1'b0;
				master0_wb_data_i <= ~32'b0;
			end
			
		endcase
	end

	// Master 1
	always @(*) begin
		case (1'b1)
			master1_slave0_select: begin
				master1_wb_ack_i <= master1_slave0_wb_ack_i;
				master1_wb_stall_i <= master1_slave0_wb_stall_i;
				master1_wb_error_i <= master1_slave0_wb_error_i;
				master1_wb_data_i <= master1_slave0_wb_data_i;
			end
			
			master1_slave1_select: begin
				master1_wb_ack_i <= master1_slave1_wb_ack_i;
				master1_wb_stall_i <= master1_slave1_wb_stall_i;
				master1_wb_error_i <= master1_slave1_wb_error_i;
				master1_wb_data_i <= master1_slave1_wb_data_i;
			end
			
			master1_slave2_select: begin
				master1_wb_ack_i <= master1_slave2_wb_ack_i;
				master1_wb_stall_i <= master1_slave2_wb_stall_i;
				master1_wb_error_i <= master1_slave2_wb_error_i;
				master1_wb_data_i <= master1_slave2_wb_data_i;
			end
			
			master1_slave3_select: begin
				master1_wb_ack_i <= master1_slave3_wb_ack_i;
				master1_wb_stall_i <= master1_slave3_wb_stall_i;
				master1_wb_error_i <= master1_slave3_wb_error_i;
				master1_wb_data_i <= master1_slave3_wb_data_i;
			end
			
			master1_slave4_select: begin
				master1_wb_ack_i <= master1_slave4_wb_ack_i;
				master1_wb_stall_i <= master1_slave4_wb_stall_i;
				master1_wb_error_i <= master1_slave4_wb_error_i;
				master1_wb_data_i <= master1_slave4_wb_data_i;
			end
			
			default: begin
				master1_wb_ack_i <= master1_wb_cyc_o;
				master1_wb_stall_i <= 1'b0;
				master1_wb_error_i <= 1'b0;
				master1_wb_data_i <= ~32'b0;
			end
			
		endcase
	end

	// Master 2
	always @(*) begin
		case (1'b1)
			master2_slave0_select: begin
				master2_wb_ack_i <= master2_slave0_wb_ack_i;
				master2_wb_stall_i <= master2_slave0_wb_stall_i;
				master2_wb_error_i <= master2_slave0_wb_error_i;
				master2_wb_data_i <= master2_slave0_wb_data_i;
			end
			
			master2_slave1_select: begin
				master2_wb_ack_i <= master2_slave1_wb_ack_i;
				master2_wb_stall_i <= master2_slave1_wb_stall_i;
				master2_wb_error_i <= master2_slave1_wb_error_i;
				master2_wb_data_i <= master2_slave1_wb_data_i;
			end
			
			master2_slave2_select: begin
				master2_wb_ack_i <= master2_slave2_wb_ack_i;
				master2_wb_stall_i <= master2_slave2_wb_stall_i;
				master2_wb_error_i <= master2_slave2_wb_error_i;
				master2_wb_data_i <= master2_slave2_wb_data_i;
			end
			
			master2_slave3_select: begin
				master2_wb_ack_i <= master2_slave3_wb_ack_i;
				master2_wb_stall_i <= master2_slave3_wb_stall_i;
				master2_wb_error_i <= master2_slave3_wb_error_i;
				master2_wb_data_i <= master2_slave3_wb_data_i;
			end
			
			master2_slave4_select: begin
				master2_wb_ack_i <= master2_slave4_wb_ack_i;
				master2_wb_stall_i <= master2_slave4_wb_stall_i;
				master2_wb_error_i <= master2_slave4_wb_error_i;
				master2_wb_data_i <= master2_slave4_wb_data_i;
			end
			
			default: begin
				master2_wb_ack_i <= master2_wb_cyc_o;
				master2_wb_stall_i <= 1'b0;
				master2_wb_error_i <= 1'b0;
				master2_wb_data_i <= ~32'b0;
			end
			
		endcase
	end

	// Master 3
	always @(*) begin
		case (1'b1)
			master3_slave0_select: begin
				master3_wb_ack_i <= master3_slave0_wb_ack_i;
				master3_wb_stall_i <= master3_slave0_wb_stall_i;
				master3_wb_error_i <= master3_slave0_wb_error_i;
				master3_wb_data_i <= master3_slave0_wb_data_i;
			end
			
			master3_slave1_select: begin
				master3_wb_ack_i <= master3_slave1_wb_ack_i;
				master3_wb_stall_i <= master3_slave1_wb_stall_i;
				master3_wb_error_i <= master3_slave1_wb_error_i;
				master3_wb_data_i <= master3_slave1_wb_data_i;
			end
			
			master3_slave2_select: begin
				master3_wb_ack_i <= master3_slave2_wb_ack_i;
				master3_wb_stall_i <= master3_slave2_wb_stall_i;
				master3_wb_error_i <= master3_slave2_wb_error_i;
				master3_wb_data_i <= master3_slave2_wb_data_i;
			end
			
			master3_slave3_select: begin
				master3_wb_ack_i <= master3_slave3_wb_ack_i;
				master3_wb_stall_i <= master3_slave3_wb_stall_i;
				master3_wb_error_i <= master3_slave3_wb_error_i;
				master3_wb_data_i <= master3_slave3_wb_data_i;
			end
			
			master3_slave4_select: begin
				master3_wb_ack_i <= master3_slave4_wb_ack_i;
				master3_wb_stall_i <= master3_slave4_wb_stall_i;
				master3_wb_error_i <= master3_slave4_wb_error_i;
				master3_wb_data_i <= master3_slave4_wb_data_i;
			end
			
			default: begin
				master3_wb_ack_i <= master3_wb_cyc_o;
				master3_wb_stall_i <= 1'b0;
				master3_wb_error_i <= 1'b0;
				master3_wb_data_i <= ~32'b0;
			end
			
		endcase
	end

	// assign probe_master0_currentSlave = master0_wb_adr_o[26:24];
	// assign probe_master1_currentSlave = master1_wb_adr_o[26:24];
	// assign probe_master2_currentSlave = master2_wb_adr_o[26:24];
	// assign probe_master3_currentSlave = master3_wb_adr_o[26:24];

	assign probe_master0_currentSlave = master0_wb_adr_o[25:24];
	assign probe_master1_currentSlave = master1_wb_adr_o[25:24];
	assign probe_master2_currentSlave = master2_wb_adr_o[25:24];
	assign probe_master3_currentSlave = master3_wb_adr_o[25:24];

endmodulemodule WishboneMultiMasterSlave (
		input wire wb_clk_i,
		input wire wb_rst_i,

		// Master 0
		input wire master0_wb_cyc_o,
		input wire master0_wb_stb_o,
		input wire master0_wb_we_o,
		input wire[3:0] master0_wb_sel_o,
		input wire[31:0] master0_wb_data_o,
		input wire[23:0] master0_wb_adr_o,
		output wire master0_wb_ack_i,
		output wire master0_wb_stall_i,
		output wire master0_wb_error_i,
		output wire[31:0] master0_wb_data_i,

		// Master 1
		input wire master1_wb_cyc_o,
		input wire master1_wb_stb_o,
		input wire master1_wb_we_o,
		input wire[3:0] master1_wb_sel_o,
		input wire[31:0] master1_wb_data_o,
		input wire[23:0] master1_wb_adr_o,
		output wire master1_wb_ack_i,
		output wire master1_wb_stall_i,
		output wire master1_wb_error_i,
		output wire[31:0] master1_wb_data_i,

		// Master 2
		input wire master2_wb_cyc_o,
		input wire master2_wb_stb_o,
		input wire master2_wb_we_o,
		input wire[3:0] master2_wb_sel_o,
		input wire[31:0] master2_wb_data_o,
		input wire[23:0] master2_wb_adr_o,
		output wire master2_wb_ack_i,
		output wire master2_wb_stall_i,
		output wire master2_wb_error_i,
		output wire[31:0] master2_wb_data_i,

		// Master 3
		input wire master3_wb_cyc_o,
		input wire master3_wb_stb_o,
		input wire master3_wb_we_o,
		input wire[3:0] master3_wb_sel_o,
		input wire[31:0] master3_wb_data_o,
		input wire[23:0] master3_wb_adr_o,
		output wire master3_wb_ack_i,
		output wire master3_wb_stall_i,
		output wire master3_wb_error_i,
		output wire[31:0] master3_wb_data_i,

		// Slave
		output wire slave_cyc_i,
		output wire slave_stb_i,
		output wire slave_we_i,
		output wire[3:0] slave_sel_i,
		output wire[31:0] slave_data_i,
		output wire[23:0] slave_adr_i,
		input wire slave_ack_o,
		input wire slave_stall_o,
		input wire slave_error_o,
		input wire[31:0] slave_data_o,

		output wire[1:0] probe_currentMaster
	);

	wire[1:0] currentMaster;
	MasterArbiter arbiter(
		.clk(wb_clk_i),
		.rst(wb_rst_i),
		.request({ master3_wb_cyc_o, master2_wb_cyc_o, master1_wb_cyc_o, master0_wb_cyc_o }),
		.masterSelected(currentMaster));
	
	wire master0Select = currentMaster == 2'h0;
	wire master1Select = currentMaster == 2'h1;
	wire master2Select = currentMaster == 2'h2;
	wire master3Select = currentMaster == 2'h3;
	
	assign slave_cyc_i =  master1Select ? master1_wb_cyc_o : 
						  master2Select ? master2_wb_cyc_o : 
						  master3Select ? master3_wb_cyc_o :
							  			  master0_wb_cyc_o;
	assign slave_stb_i =  master1Select ? master1_wb_stb_o : 
						  master2Select ? master2_wb_stb_o : 
						  master3Select ? master3_wb_stb_o :
							  			  master0_wb_stb_o;
	assign slave_we_i =   master1Select ? master1_wb_we_o : 
						  master2Select ? master2_wb_we_o : 
						  master3Select ? master3_wb_we_o :
							  			  master0_wb_we_o;
	assign slave_sel_i =  master1Select ? master1_wb_sel_o : 
						  master2Select ? master2_wb_sel_o : 
						  master3Select ? master3_wb_sel_o :
							  			  master0_wb_sel_o;
	assign slave_data_i = master1Select ? master1_wb_data_o : 
						  master2Select ? master2_wb_data_o : 
						  master3Select ? master3_wb_data_o :
							  			  master0_wb_data_o;
	assign slave_adr_i =  master1Select ? master1_wb_adr_o : 
						  master2Select ? master2_wb_adr_o : 
						  master3Select ? master3_wb_adr_o :
							  			  master0_wb_adr_o;

	// Master 0
	assign master0_wb_ack_i   = slave_ack_o;
	assign master0_wb_stall_i = slave_stall_o;
	assign master0_wb_error_i = slave_error_o;
	assign master0_wb_data_i  = slave_data_o;

	// Master 1
	assign master1_wb_ack_i   = slave_ack_o;
	assign master1_wb_stall_i = slave_stall_o;
	assign master1_wb_error_i = slave_error_o;
	assign master1_wb_data_i  = slave_data_o;

	// Master 2
	assign master2_wb_ack_i   = slave_ack_o;
	assign master2_wb_stall_i = slave_stall_o;
	assign master2_wb_error_i = slave_error_o;
	assign master2_wb_data_i  = slave_data_o;

	// Master 3
	assign master3_wb_ack_i   = slave_ack_o;
	assign master3_wb_stall_i = slave_stall_o;
	assign master3_wb_error_i = slave_error_o;
	assign master3_wb_data_i  = slave_data_o;

	// Assign logic probes
	assign probe_currentMaster = currentMaster;
endmodulemodule MasterArbiter (
		input wire clk,
		input wire rst,

		input wire[3:0] request,
		output wire[1:0] masterSelected
	);

	localparam MASTER0 = 2'h0;
	localparam MASTER1 = 2'h1;
	localparam MASTER2 = 2'h2;
	localparam MASTER3 = 2'h3;

	reg[1:0] currentMaster = MASTER0;
	reg[1:0] nextMaster;

	always @(*) begin
		nextMaster = currentMaster;

		case (currentMaster)
			MASTER0: begin
				if (!request[0]) begin
					if (request[1]) nextMaster = MASTER1;
					else if (request[2]) nextMaster = MASTER2;
					else if (request[3]) nextMaster = MASTER3;
				end
			end

			MASTER1: begin
				if (!request[1]) begin
					if (request[2]) nextMaster = MASTER2;
					else if (request[3]) nextMaster = MASTER3;
					else if (request[0]) nextMaster = MASTER0;
				end
			end

			MASTER2: begin
				if (!request[2]) begin
					if (request[3]) nextMaster = MASTER3;
					else if (request[0]) nextMaster = MASTER0;
					else if (request[1]) nextMaster = MASTER1;
				end
			end

			MASTER3: begin
				if (!request[3]) begin
					if (request[0]) nextMaster = MASTER0;
					else if (request[1]) nextMaster = MASTER1;
					else if (request[2]) nextMaster = MASTER2;
				end
			end
		endcase
	end

	always @(posedge clk) begin
		if (rst) currentMaster <= MASTER0;
		else currentMaster <= nextMaster;
	end

	assign masterSelected = nextMaster;

endmodulemodule FIFO
	#(
		parameter WORD_SIZE = 8,
		parameter BUFFER_SIZE = 256	// If this is not a power of two, the actual buffer size will be the smallest power of two greater than BUFFER_SIZE
	)(
		input wire clk,
		input wire rst,
		input wire [WORD_SIZE-1:0] dataIn,
		input wire we,

		output wire [WORD_SIZE-1:0] dataOut,
		input wire oe,
		
		output wire isData,
		output wire bufferFull,
		output wire dataLost
    );

	localparam ADDRESS_SIZE = $clog2(BUFFER_SIZE);
	localparam DEPTH = 1 << ADDRESS_SIZE;

	reg we_buffered = 1'b0;
	reg oe_buffered = 1'b0;
	reg[WORD_SIZE-1:0] dataIn_buffered = {WORD_SIZE{1'b0}};
	reg[WORD_SIZE-1:0] dataOut_buffered;

	reg[ADDRESS_SIZE-1:0] startPointer = {ADDRESS_SIZE{1'b0}};
	reg[ADDRESS_SIZE-1:0] endPointer = {ADDRESS_SIZE{1'b0}};
	reg[WORD_SIZE-1:0] buffer [0:DEPTH-1];

	wire[ADDRESS_SIZE-1:0] nextStartPointer = startPointer + 1;
	wire[ADDRESS_SIZE-1:0] nextEndPointer = endPointer + 1;

	reg lastWriteLostData = 1'b0;


	always @(posedge clk) begin
		if (rst) begin
			we_buffered <= 1'b0;
			oe_buffered <= 1'b0;
			dataIn_buffered <= {WORD_SIZE{1'b0}};
		end else begin
			we_buffered <= we;
			oe_buffered <= oe;
			dataIn_buffered <= dataIn;
		end
	end

	always @(negedge clk) begin
		if (rst) begin
			startPointer <= {ADDRESS_SIZE{1'b0}};
			endPointer <= {ADDRESS_SIZE{1'b0}};
			lastWriteLostData <= 1'b0;
			dataOut_buffered <= {WORD_SIZE{1'b0}};
		end else begin
			if (oe_buffered) begin
				if (isData) begin
					startPointer <= nextStartPointer;
					dataOut_buffered <= buffer[nextStartPointer];
				end else begin
					dataOut_buffered <= {WORD_SIZE{1'b0}};
				end
			end

			if (we_buffered) begin
				// TODO: Should we allow the buffer to overwrite itself when a write occurs and it is already full
				if (!bufferFull) begin
					buffer[endPointer] <= dataIn_buffered;					
					endPointer <= nextEndPointer;
					lastWriteLostData <= 1'b0;

					if (!isData) dataOut_buffered <= dataIn_buffered;
				end else begin
					lastWriteLostData <= 1'b1;
				end
			end
		end
	end

	assign dataOut = dataOut_buffered;

	assign isData = startPointer != endPointer;
	assign bufferFull = nextEndPointer == startPointer;
	assign dataLost = lastWriteLostData;	

endmodule
module Mux #(
		parameter WIDTH = 1,
		parameter INPUTS = 2,
		parameter DEFAULT = 'b0
	)(
		input wire[INPUTS-1:0] select,
		input wire[(WIDTH*INPUTS)-1:0] in,
		output reg[WIDTH-1:0] out,
		output wire outputEnable
	);
	
	generate
		if (INPUTS == 1) begin
			always @(*) begin
				case (1'b1)
					select[0]: out <= in[WIDTH-1:0];
					default: out <= DEFAULT;
				endcase
			end
		end else if (INPUTS == 2) begin
			always @(*) begin
				case (1'b1)
					select[0]: out <= in[WIDTH-1:0];
					select[1]: out <= in[(1 * WIDTH) + WIDTH - 1:1 * WIDTH];
					default: out <= DEFAULT;
				endcase
			end
		end else if (INPUTS == 3) begin
			always @(*) begin
				case (1'b1)
					select[0]: out <= in[WIDTH-1:0];
					select[1]: out <= in[(1 * WIDTH) + WIDTH - 1:1 * WIDTH];
					select[2]: out <= in[(2 * WIDTH) + WIDTH - 1:2 * WIDTH];
					default: out <= DEFAULT;
				endcase
			end
		end else if (INPUTS == 4) begin
			always @(*) begin
				case (1'b1)
					select[0]: out <= in[WIDTH-1:0];
					select[1]: out <= in[(1 * WIDTH) + WIDTH - 1:1 * WIDTH];
					select[2]: out <= in[(2 * WIDTH) + WIDTH - 1:2 * WIDTH];
					select[3]: out <= in[(3 * WIDTH) + WIDTH - 1:3 * WIDTH];
					default: out <= DEFAULT;
				endcase
			end
		end else if (INPUTS == 5) begin
			always @(*) begin
				case (1'b1)
					select[0]: out <= in[WIDTH-1:0];
					select[1]: out <= in[(1 * WIDTH) + WIDTH - 1:1 * WIDTH];
					select[2]: out <= in[(2 * WIDTH) + WIDTH - 1:2 * WIDTH];
					select[3]: out <= in[(3 * WIDTH) + WIDTH - 1:3 * WIDTH];
					select[4]: out <= in[(4 * WIDTH) + WIDTH - 1:4 * WIDTH];
					default: out <= DEFAULT;
				endcase
			end
		end else if (INPUTS == 6) begin
			always @(*) begin
				case (1'b1)
					select[0]: out <= in[WIDTH-1:0];
					select[1]: out <= in[(1 * WIDTH) + WIDTH - 1:1 * WIDTH];
					select[2]: out <= in[(2 * WIDTH) + WIDTH - 1:2 * WIDTH];
					select[3]: out <= in[(3 * WIDTH) + WIDTH - 1:3 * WIDTH];
					select[4]: out <= in[(4 * WIDTH) + WIDTH - 1:4 * WIDTH];
					select[5]: out <= in[(5 * WIDTH) + WIDTH - 1:5 * WIDTH];
					default: out <= DEFAULT;
				endcase
			end
		end else if (INPUTS == 7) begin
			always @(*) begin
				case (1'b1)
					select[0]: out <= in[WIDTH-1:0];
					select[1]: out <= in[(1 * WIDTH) + WIDTH - 1:1 * WIDTH];
					select[2]: out <= in[(2 * WIDTH) + WIDTH - 1:2 * WIDTH];
					select[3]: out <= in[(3 * WIDTH) + WIDTH - 1:3 * WIDTH];
					select[4]: out <= in[(4 * WIDTH) + WIDTH - 1:4 * WIDTH];
					select[5]: out <= in[(5 * WIDTH) + WIDTH - 1:5 * WIDTH];
					select[6]: out <= in[(6 * WIDTH) + WIDTH - 1:6 * WIDTH];
					default: out <= DEFAULT;
				endcase
			end
		end else if (INPUTS == 8) begin
			always @(*) begin
				case (1'b1)
					select[0]: out <= in[WIDTH-1:0];
					select[1]: out <= in[(1 * WIDTH) + WIDTH - 1:1 * WIDTH];
					select[2]: out <= in[(2 * WIDTH) + WIDTH - 1:2 * WIDTH];
					select[3]: out <= in[(3 * WIDTH) + WIDTH - 1:3 * WIDTH];
					select[4]: out <= in[(4 * WIDTH) + WIDTH - 1:4 * WIDTH];
					select[5]: out <= in[(5 * WIDTH) + WIDTH - 1:5 * WIDTH];
					select[6]: out <= in[(6 * WIDTH) + WIDTH - 1:6 * WIDTH];
					select[7]: out <= in[(7 * WIDTH) + WIDTH - 1:7 * WIDTH];
					default: out <= DEFAULT;
				endcase
			end
		end else begin
			// integer i;
			// always @(*) begin
			// 	for (i = 0; i < INPUTS; i = i + 1) begin
			// 		if (select[i]) out <= in[(i * WIDTH) + WIDTH - 1:i * WIDTH];
			// 	end
			// end
		end
	endgenerate

	assign outputEnable = |select;

endmodulemodule ShiftRegister #(
		parameter WIDTH = 8
	)(
		input wire clk,
		input wire rst,

		input wire loadEnable,
		input wire shiftInEnable,
		input wire shiftOutEnable,
		input wire msbFirst,

		input  wire[WIDTH-1:0] parallelIn,
		output wire[WIDTH-1:0] parallelOut,
		input  wire serialIn,
		output wire serialOut
	);

	reg[WIDTH-1:0] data;
	reg outputBit = 1'b0;
	wire[WIDTH-1:0] nextData;

	generate
		if (WIDTH == 1) begin
			assign nextData = serialIn;
		end else begin
			assign nextData = msbFirst ? { data[WIDTH-2:0], serialIn } : { serialIn, data[WIDTH-1:1] };
		end
	endgenerate
	

	always @(posedge clk) begin
		if (rst) begin
			data <= {WIDTH{1'b0}};
			outputBit <= 1'b0;
		end else if (loadEnable) begin
			data <= parallelIn;
			outputBit <= msbFirst ? parallelIn[WIDTH-1] : parallelIn[0];
		end	else if (shiftInEnable) begin
			data <= nextData;
			if (shiftOutEnable) outputBit <= msbFirst ? nextData[WIDTH-1] : nextData[0];
		end else if (shiftOutEnable) outputBit <= msbFirst ? data[WIDTH-1] : data[0];

	end
		
	assign parallelOut = data;
	assign serialOut = outputBit;

endmodulemodule Counter #(
		parameter WIDTH = 8, 	// Width of the output
		parameter DIV = 0, 		// number of bits to use as divisor
		parameter TOP = 0, 		// max value, 0 = none		
		parameter UP = 1 		// direction to count, use 1 for up and 0 for down
	)(
		input wire clk,
		input wire rst,
		input wire halt,
		output reg [WIDTH-1:0] value
	);
  
	reg [WIDTH + DIV - 1:0] counter = 'b0;

	always @(posedge clk) begin		
		if (TOP != 'b0) begin
			if (rst || (counter[WIDTH + DIV - 1:DIV] == TOP)) counter = 'b0;
			else begin
				if (!halt) begin
					if (UP) counter = counter + 1;
					else counter = counter - 1;
				end
			end
		end else begin
			if (rst) begin
				counter = 'b0;
			end else begin
				if (!halt) begin
					if (UP) counter = counter + 1;
					else counter = counter - 1;
				end
			end
		end
		
		value = counter[WIDTH + DIV - 1:DIV];
	end

endmodule
(* blackbox *)
module Art (

		inout vccd1,	// User area 1 1.8V supply
		inout vssd1//,	// User area 1 digital ground

		//output wire dumyPin
	);
	
endmodule`default_nettype none

`timescale 1 ns / 1 ps

















































































































//`define RV32I_NOP 32'h00000013

`timescale 1 ns / 1 ps





































































































































module UserSpace(
		input wire clk,
		input wire rst,

		input wire [127:0] la_data_in_user,
		output wire [127:0] la_data_out_user,
		input wire [127:0] la_oenb_user,

		output wire [(19 + 19)-1:0] user_io_oeb,
		input wire [(19 + 19)-1:0] user_io_in,
		output wire [(19 + 19)-1:0] user_io_out,
		inout wire [(19 + 19)-10:0] mprj_analog_io,

		output wire[2:0] user_irq_core,

		input wire[31:0] wbAddress,
		input wire[3:0] wbByteSelect,
		input wire wbEnable,
		input wire wbWriteEnable,
		input wire[31:0] wbDataWrite,
		output wire[31:0] wbDataRead,
		output wire wbBusy,

		input wire succesOutput,
		input wire nextTestOutput
	);

	// Dispaly message with result of each test, ending the simulation if a test fails
	reg[31:0] testCounter = 0;
	always @(succesOutput, nextTestOutput) begin
		#1
		if (nextTestOutput) begin
			if (succesOutput) begin
				$display("%c[1;92mPassed test: %d%c[0m", 27, testCounter, 27);
			end	else begin
				$display("%c[1;31mFailed test: %d%c[0m", 27, testCounter, 27);
				#500
				$finish;
			end
			testCounter <= testCounter + 1;
		end
	end

	reg power1, power2;
	reg power3, power4;

	initial begin		// Power-up sequence
		power1 <= 1'b0;
		power2 <= 1'b0;
		power3 <= 1'b0;
		power4 <= 1'b0;
		#100;
		power1 <= 1'b1;
		#100;
		power2 <= 1'b1;
		#100;
		power3 <= 1'b1;
		#100;	
		power4 <= 1'b1;
	end

	wire VDD3V3;
	wire VDD1V8;
	wire VSS;
	
	assign VDD3V3 = power1;
	assign VDD1V8 = power2;
	assign VSS = 1'b0;

	 // Exported Wishbone Bus (user area facing)
	wire 	mprj_cyc_o_user;
	wire 	mprj_stb_o_user;
	wire 	mprj_we_o_user;
	wire [3:0]  mprj_sel_o_user;
	wire [31:0] mprj_adr_o_user;
	wire [31:0] mprj_dat_o_user;
	wire [31:0] mprj_dat_i_user;
	wire	mprj_ack_i_user;
	
	Core_WBInterface #(.ADDRESS_WIDTH(32)) mprj_wb_interface (
		// Wishbone master interface
		.wb_clk_i(clk),
		.wb_rst_i(rst),
		.wb_cyc_o(mprj_cyc_o_user),
		.wb_stb_o(mprj_stb_o_user),
		.wb_we_o(mprj_we_o_user),
		.wb_sel_o(mprj_sel_o_user),
		.wb_data_o(mprj_dat_o_user),
		.wb_adr_o(mprj_adr_o_user),
		.wb_ack_i(mprj_ack_i_user),
		.wb_stall_i(1'b0),
		.wb_error_i(1'b0),
		.wb_data_i(mprj_dat_i_user),

		// Memory interface from core
		.wbAddress(wbAddress),
		.wbByteSelect(wbByteSelect),
		.wbEnable(wbEnable),
		.wbWriteEnable(wbWriteEnable),
		.wbDataWrite(wbDataWrite),
		.wbDataRead(wbDataRead),
		.wbBusy(wbBusy)
	);

	user_project_wrapper mprj ( 
		.vdda1(VDD3V3),		// User area 1 3.3V power
		.vdda2(VDD3V3),		// User area 2 3.3V power
		.vssa1(VSS),		// User area 1 analog ground
		.vssa2(VSS),		// User area 2 analog ground
		.vccd1(VDD1V8),		// User area 1 1.8V power
		.vccd2(VDD1V8),		// User area 2 1.8V power
		.vssd1(VSS),		// User area 1 digital ground
		.vssd2(VSS),		// User area 2 digital ground

		.wb_clk_i(clk),
		.wb_rst_i(rst),

		// Management SoC Wishbone bus (exported)
		.wbs_cyc_i(mprj_cyc_o_user),
		.wbs_stb_i(mprj_stb_o_user),
		.wbs_we_i(mprj_we_o_user),
		.wbs_sel_i(mprj_sel_o_user),
		.wbs_adr_i(mprj_adr_o_user),
		.wbs_dat_i(mprj_dat_o_user),
		.wbs_ack_o(mprj_ack_i_user),
		.wbs_dat_o(mprj_dat_i_user),

		// GPIO pad 3-pin interface (plus analog)
		.io_in (user_io_in),
		.io_out(user_io_out),
		.io_oeb(user_io_oeb),
		.analog_io(mprj_analog_io),

		// Logic analyzer
		.la_data_in(la_data_in_user),
		.la_data_out(la_data_out_user),
		.la_oenb(la_oenb_user),

		// Independent clock
		.user_clock2(clk),

		// IRQ
		.user_irq(user_irq_core)
	);

endmodule

module userSpace_tb;
	reg clk;
	reg rst;

	reg [127:0] la_data_in_user = 128'b0;  // From CPU to MPRJ
	wire [127:0] la_data_out_user; // From MPRJ to CPU
	reg [127:0] la_oenb_user = ~128'b0;	 // From CPU to MPRJ

	wire [(19 + 19)-1:0] user_io_oeb;
	reg [(19 + 19)-1:0] user_io_in = 'b0;
	wire [(19 + 19)-1:0] user_io_out;
	wire [(19 + 19)-10:0] mprj_analog_io;

	reg[31:0] wbAddress = 32'b0;
	reg[3:0] wbByteSelect = 4'b0;
	reg wbEnable = 1'b0;
	reg wbWriteEnable = 1'b0;
	reg[31:0] wbDataWrite = 32'b0;
	wire[31:0] wbDataRead;
	wire wbBusy;

	reg succesOutput = 1'b1;
	reg nextTestOutput = 1'b0;

	wire [2:0]   user_irq_core;

	initial begin
		$dumpfile("userSpace.vcd");
		$dumpvars(0, userSpace_tb);
		
	repeat (100) begin
		repeat (1000) @(posedge clk);
	end
	$display("%c[1;35m",27);
	


		$display ("Monitor: Timeout, Core PC Test (RTL) Failed");
	
	$display("%c[0m",27);

		$finish;
	end

	reg[6:0] tmp;
	reg[31:0] testValue = 32'b0;
	reg[31:0] initialInstructionCount = 32'b0;
	initial begin
		@(negedge rst);
		#100

		// Run tests
		// Setup test data in sram and make sure the test data has been written correctly
		// If it isn't probably run a specific memory test, rather than this one
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30000000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30000000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= { ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 };
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30000000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30000000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h30000000) + {(32'h40), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h30000000) + {(32'h40), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= { ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 };
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h30000000) + {(32'h40), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h30000000) + {(32'h40), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h30000000) + {(32'h41), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h30000000) + {(32'h41), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= { ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 };
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h30000000) + {(32'h41), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h30000000) + {(32'h41), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h30000000) + {(32'h42), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h30000000) + {(32'h42), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= { ((-32'h4) >> (20)) & 32'h1, ((-32'h4) >> (1)) & ((32'h1 << (10 - 1 + 1)) - 32'h1), ((-32'h4) >> (11)) & 32'h1, ((-32'h4) >> (12)) & ((32'h1 << (19 - 12 + 1)) - 32'h1), 5'h00, 7'b1101111 };
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h30000000) + {(32'h42), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h30000000) + {(32'h42), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((-32'h4) >> (20)) & 32'h1, ((-32'h4) >> (1)) & ((32'h1 << (10 - 1 + 1)) - 32'h1), ((-32'h4) >> (11)) & 32'h1, ((-32'h4) >> (12)) & ((32'h1 << (19 - 12 + 1)) - 32'h1), 5'h00, 7'b1101111 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;
		

		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31000000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31000000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= { ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 };
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31000000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31000000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h31000000) + {(32'h40), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h31000000) + {(32'h40), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= { ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 };
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h31000000) + {(32'h40), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h31000000) + {(32'h40), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h31000000) + {(32'h41), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h31000000) + {(32'h41), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= { ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 };
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h31000000) + {(32'h41), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h31000000) + {(32'h41), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h31000000) + {(32'h42), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h31000000) + {(32'h42), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= { ((-32'h4) >> (20)) & 32'h1, ((-32'h4) >> (1)) & ((32'h1 << (10 - 1 + 1)) - 32'h1), ((-32'h4) >> (11)) & 32'h1, ((-32'h4) >> (12)) & ((32'h1 << (19 - 12 + 1)) - 32'h1), 5'h00, 7'b1101111 };
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h31000000) + {(32'h42), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h31000000) + {(32'h42), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((-32'h4) >> (20)) & 32'h1, ((-32'h4) >> (1)) & ((32'h1 << (10 - 1 + 1)) - 32'h1), ((-32'h4) >> (11)) & 32'h1, ((-32'h4) >> (12)) & ((32'h1 << (19 - 12 + 1)) - 32'h1), 5'h00, 7'b1101111 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Test core 0
		// Read that the config defaulted to 0
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h0));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Read that the program counter defaulted to 0x0000_0000
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30810000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30810000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h0));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Step PC
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30810008) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30810008) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);

		// Read that the PC stepped once
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30810000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30810000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h4));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Check that a NOP was read
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30810010) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30810010) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Jump PC
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30810004) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30810004) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h100;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);

		// Read that the PC jumped correctly
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30810000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30810000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h104));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Let the core run
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h1;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
		#200
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);

		// Make sure the core halted
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h0));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Check that the core has run
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h30818000) + {(30'hC02), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h30818000) + {(30'hC02), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	initialInstructionCount <= wbDataRead;
		
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (initialInstructionCount > 1 && initialInstructionCount != ~32'h0);
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Let the core run
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h1;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
		#200
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);

		// Make sure the core halted
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h0));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Check that the core has been restarted
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h30818000) + {(30'hC02), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h30818000) + {(30'hC02), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
		
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue > initialInstructionCount);
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Check that the PC has increased should be either 0x104 or 0x108
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h30810000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h30810000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
		
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == 32'h104 || testValue == 32'h108);
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Test core 1
		// Read that the config defaulted to 0
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h0));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Read that the program counter defaulted to 0x0000_0000
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31810000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31810000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h0));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Step PC
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31810008) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31810008) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);

		// Read that the PC stepped once
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31810000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31810000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h4));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Check that an NOP was read
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31810010) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31810010) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == ({ ((32'h0) >> (0)) & ((32'h1 << (11 - 0 + 1)) - 32'h1), 5'h00, 3'b000, 5'h00, 7'b0010011 }));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Jump PC
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31810004) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31810004) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h100;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);

		// Read that the PC jumped correctly
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31810000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31810000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h104));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Let the core run
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h1;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
		#200
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);

		// Make sure the core halted
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h0));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Check that the core is running
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h31818000) + {(30'hC02), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h31818000) + {(30'hC02), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	initialInstructionCount <= wbDataRead;
		
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (initialInstructionCount > 1 && initialInstructionCount != ~32'h0);
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		// Let the core run
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h1;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
		#200
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= 32'h0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);

		// Make sure the core halted
		
	
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31800000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31800000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
	
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == (32'h0));
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;


		// Check that the core has been restarted
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= ((32'h31818000) + {(30'hC02), 2'b00}) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= (((32'h31818000) + {(30'hC02), 2'b00}) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
		
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue > initialInstructionCount);
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;
		
		// Check that the PC has increased should be either 0x104 or 0x108
		
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= 32'h30000000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b1;
	wbDataWrite <= (32'h31810000) & 32'hFFFF8000;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	
	@(negedge clk)
	#1
	wait(!wbBusy);
	wbAddress <= ((32'h31810000) & 32'h00007FFF) | 32'h30008000;
	wbByteSelect <= 4'b1111;
	wbWriteEnable <= 1'b0;
	wbEnable <= 1'b1;
	@(posedge clk)
	@(posedge clk)
	@(posedge clk)
	wait(!wbBusy);
	testValue <= wbDataRead;
		
	@(negedge clk)
	#1
	if (succesOutput) succesOutput <= (testValue == 32'h104 || testValue == 32'h108);
	nextTestOutput <= 1'b1;
	@(posedge clk);
	@(negedge clk);
	nextTestOutput <= 1'b0;

		
	#100
	if (succesOutput) begin
		$display("%c[1;92m",27);
		


			$display("Monitor: Core PC Test (RTL) Passed");
		
		$display("%c[0m",27);
	end else begin
		$display("%c[1;31m",27);
		


			$display ("Monitor: Core PC Test (RTL) Failed");
		
		$display("%c[0m",27);
	end
	    $finish;
	end

	// External clock is used by default.  Make this artificially fast for the
	// simulation.  Normally this would be a slow clock and the digital PLL
	// would be the fast clock.
	always #12.5 clk <= (clk === 1'b0);

	initial begin
		rst <= 1'b1;
		#2000;
		rst <= 1'b0; // Release reset
	end

	UserSpace userSpace(
		.clk(clk),
		.rst(rst),
		.la_data_in_user(la_data_in_user),
		.la_data_out_user(la_data_out_user),
		.la_oenb_user(la_oenb_user),
		.user_io_oeb(user_io_oeb),
		.user_io_in(user_io_in),
		.user_io_out(user_io_out),
		.mprj_analog_io(mprj_analog_io),
		.user_irq_core(user_irq_core),
		.wbAddress(wbAddress),
		.wbByteSelect(wbByteSelect),
		.wbEnable(wbEnable),
		.wbWriteEnable(wbWriteEnable),
		.wbDataWrite(wbDataWrite),
		.wbDataRead(wbDataRead),
		.wbBusy(wbBusy),
		.succesOutput(succesOutput),
		.nextTestOutput(nextTestOutput));

endmodule
`default_nettype wire
